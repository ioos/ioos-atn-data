netcdf NCEI_test.3 {
dimensions:
	obs = 5217 ;
variables:
	int crs ;
		crs:epsg_code = "EPSG:4326" ;
		crs:grid_mapping_name = "latitude_longitude" ;
		crs:inverse_flattening = 298.257223563 ;
		crs:ioos_category = "Other" ;
		crs:long_name = "http://www.opengis.net/def/crs/EPSG/0/4326" ;
		crs:semi_major_axis = 6378137. ;
	double ellipse_orientation(obs) ;
		ellipse_orientation:_FillValue = -9999.9 ;
		ellipse_orientation:coordinates = "time z lon lat" ;
		ellipse_orientation:long_name = "Platform identifier" ;
		ellipse_orientation:units = "degrees" ;
		ellipse_orientation:comment = "The angle in degrees of the ellipse from true north, proceeding clockwise (0 to 360). A blank field represents 0 degrees." ;
		ellipse_orientation:instrument = "instrument_location" ;
		ellipse_orientation:platform = "platform" ;
	double error_radius(obs) ;
		error_radius:_FillValue = -9999.9 ;
		error_radius:coordinates = "time z lon lat" ;
		error_radius:long_name = "Error radius" ;
		error_radius:units = "m" ;
		error_radius:comment = "If the position is best represented as a circle, this field gives the radius of that circle in meters." ;
		error_radius:instrument = "instrument_location" ;
		error_radius:platform = "platform" ;
	string instrument_location ;
		instrument_location:long_name = "Wildlife Computers Splash 10" ;
		instrument_location:location_type = "argos / modeled" ;
		instrument_location:comment = "Location" ;
		instrument_location:manufacturer = "Wildlife Computers" ;
		instrument_location:make_model = "Splash 10" ;
		instrument_location:calibration_date = "" ;
		instrument_location:serial_number = "18A0360" ;
	string instrument_pressure ;
		instrument_pressure:long_name = "some pressure sensor" ;
		instrument_pressure:comment = "hypothetical WC pressure sensos" ;
		instrument_pressure:manufacturer = "Wildlife Computers" ;
		instrument_pressure:make_model = "WC pressure sensor" ;
		instrument_pressure:calibration_date = "" ;
		instrument_pressure:serial_number = "XXX55544XO" ;
	string instrument_tag ;
		instrument_tag:long_name = "instrument" ;
		instrument_tag:comment = "Test comment" ;
		instrument_tag:manufacturer = "Wildlife Computers" ;
		instrument_tag:make_model = "Splash 10" ;
		instrument_tag:calibration_date = "" ;
		instrument_tag:serial_number = "18A0360" ;
	double lat(obs) ;
		lat:_FillValue = -9999.9 ;
		lat:axis = "Y" ;
		lat:_CoordinateAxisType = "Lat" ;
		lat:ioos_category = "Location" ;
		lat:long_name = "Profile Location" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:valid_max = 90. ;
		lat:valid_min = -90. ;
		lat:actual_min = 50.6209 ;
		lat:actual_max = 66.8307 ;
		lat:instrument = "instrument_location" ;
		lat:platform = "platform" ;
	string location_class(obs) ;
		location_class:coordinates = "time z lon lat" ;
		location_class:long_name = "Location Quality Code" ;
		location_class:standard_name = "quality_code" ;
		location_class:ioos_category = "Quality" ;
		location_class:comment = "Quality codes from the ARGOS satellite (in meters): G,3,2,1,0,A,B,Z. See http://www.argos-system.org/manual/3-location/34_location_classes.htm" ;
		location_class:instrument = "instrument_location" ;
		location_class:platform = "platform" ;
	double lon(obs) ;
		lon:_FillValue = -9999.9 ;
		lon:axis = "X" ;
		lon:_CoordinateAxisType = "Lon" ;
		lon:ioos_category = "Location" ;
		lon:long_name = "Profile Location" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:valid_max = 180. ;
		lon:valid_min = -180. ;
		lon:actual_min = -154.258 ;
		lon:actual_max = 160.9647 ;
		lon:instrument = "instrument_location" ;
		lon:platform = "platform" ;
	double offset(obs) ;
		offset:_FillValue = -9999.9 ;
		offset:coordinates = "time z lon lat" ;
		offset:long_name = "Offset" ;
		offset:units = "m" ;
		offset:comment = "This field is non-zero if the circle or ellipse are not centered on the (Latitude, Longitude) values on this row. \"Offset\" gives the distance in meters from (Latitude, Longitude) to the center of the ellipse." ;
	double offset_orientation(obs) ;
		offset_orientation:_FillValue = -9999.9 ;
		offset_orientation:coordinates = "time z lon lat" ;
		offset_orientation:long_name = "Offset orientation" ;
		offset_orientation:units = "degrees" ;
		offset_orientation:comment = "If the \"Offset\" field is non-zero, this field is the angle in degrees from (Latitude, Longitude) to the center of the ellipse. Zero degrees is true north; a blank field represents 0 degrees." ;
	string platform ;
		platform:cf_role = "5deb0b1d6321be14905284b8" ;
		platform:long_name = "SSL2019788KOD" ;
		platform:platform_type = "animal" ;
		platform:platform_vocabulary = "https://mmisw.org/ont/ioos/platform" ;
		platform:valid_name = "Eumetopias jubatus" ;
		platform:AphiaID = 254999LL ;
		platform:scientificname = "Eumetopias jubatus" ;
		platform:authority = "(Schreber, 1776)" ;
		platform:kingdom = "Animalia" ;
		platform:phylum = "Chordata" ;
		platform:class = "Mammalia" ;
		platform:order = "Carnivora" ;
		platform:family = "Otariidae" ;
		platform:genus = "Eumetopias" ;
		platform:taxonRankID = 220LL ;
		platform:rank = "Species" ;
		platform:superdomain = "Biota" ;
		platform:subphylum = "Vertebrata" ;
		platform:superclass = "Tetrapoda" ;
		platform:subclass = "Theria" ;
		platform:suborder = "Caniformia" ;
		platform:infraorder = "Pinnipedia" ;
		platform:species = "Eumetopias jubatus" ;
	string qartod_location_flag ;
		string qartod_location_flag:_FillValue = "0" ;
		qartod_location_flag:flag_meanings = "PASS NOT_EVALUATED SUSPECT FAIL MISSING" ;
		qartod_location_flag:flag_values = "1, 2, 3, 4, 9" ;
		qartod_location_flag:ioos_category = "Other" ;
		qartod_location_flag:long_name = "" ;
		qartod_location_flag:standard_name = "" ;
	string qartod_rollup_flag2 ;
		string qartod_rollup_flag2:_FillValue = "0" ;
		qartod_rollup_flag2:flag_meanings = "PASS NOT_EVALUATED SUSPECT FAIL MISSING" ;
		qartod_rollup_flag2:flag_values = "1, 2, 3, 4, 9" ;
		qartod_rollup_flag2:ioos_category = "Other" ;
		qartod_rollup_flag2:long_name = "" ;
		qartod_rollup_flag2:standard_name = "" ;
	string qartod_speed_flag ;
		string qartod_speed_flag:_FillValue = "0" ;
		qartod_speed_flag:flag_meanings = "PASS NOT_EVALUATED SUSPECT FAIL MISSING" ;
		qartod_speed_flag:flag_values = "1, 2, 3, 4, 9" ;
		qartod_speed_flag:ioos_category = "Other" ;
		qartod_speed_flag:long_name = "" ;
		qartod_speed_flag:standard_name = "" ;
	string qartod_time_flag ;
		string qartod_time_flag:_FillValue = "0" ;
		qartod_time_flag:flag_meanings = "PASS NOT_EVALUATED SUSPECT FAIL MISSING" ;
		qartod_time_flag:flag_values = "1, 2, 3, 4, 9" ;
		qartod_time_flag:ioos_category = "Other" ;
		qartod_time_flag:long_name = "" ;
		qartod_time_flag:standard_name = "" ;
	double semi_major_axis(obs) ;
		semi_major_axis:_FillValue = -9999.9 ;
		semi_major_axis:coordinates = "time z lon lat" ;
		semi_major_axis:long_name = "Error semi-major axis" ;
		semi_major_axis:units = "m" ;
		semi_major_axis:comment = "If the estimated position error is best expressed as an ellipse, this field gives the length in meters of the semi-major elliptical axis (one half of the major axis)." ;
		semi_major_axis:instrument = "instrument_location" ;
		semi_major_axis:platform = "platform" ;
	double semi_minor_axis(obs) ;
		semi_minor_axis:_FillValue = -9999.9 ;
		semi_minor_axis:coordinates = "time z lon lat" ;
		semi_minor_axis:long_name = "Error semi-minor axis" ;
		semi_minor_axis:units = "m" ;
		semi_minor_axis:comment = "If the estimated position error is best expressed as an ellipse, this field gives the length in meters of the semi-minor elliptical axis (one half of the minor axis)." ;
		semi_minor_axis:instrument = "instrument_location" ;
		semi_minor_axis:platform = "platform" ;
	double time(obs) ;
		time:_FillValue = -9999.9 ;
		time:units = "seconds since 1990-01-01 00:00:00Z" ;
		time:standard_name = "time" ;
		time:axis = "T" ;
		time:_CoordinateAxisType = "Time" ;
		time:calendar = "standard" ;
		time:ioos_category = "Time" ;
		time:long_name = "Time" ;
		time:actual_min = "2019-11-29T15:05:02Z" ;
		time:actual_max = "2020-04-27T08:29:22Z" ;
	int z(obs) ;
		z:_FillValue = -9999 ;
		z:axis = "Z" ;
		z:long_name = "depth" ;
		z:positive = "down" ;
		z:standard_name = "depth" ;
		z:units = "m" ;
		z:actual_min = 0. ;
		z:actual_max = 0. ;
		z:instrument = "instrument_location" ;
		z:platform = "platform" ;

// global attributes:
		:date_created = "2020-04-27T16:04:41Z" ;
		:featureType = "trajectory" ;
		:cdm_data_type = "Trajectory" ;
		:geospatial_bounds_vertical_crs = "EPSG:4326" ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_vertical_positive = "down" ;
		:naming_authority = "gov.noaa.ioos.atn" ;
		:publisher_email = "atndata@ioos.us" ;
		:publisher_name = "IOOS ATN" ;
		:publisher_url = "https://atn.ioos.us" ;
		:source = "Service Argos" ;
		:standard_name_vocabulary = "CF-v58" ;
		:geospatial_bbox = "POLYGON ((250.83 50.6209, 250.83 66.83069999999999, 159.0115000000001 66.83069999999999, 159.0115000000001 50.6209, 250.83 50.6209))" ;
		:geospatial_bounds = "POLYGON ((159.0115000000001 50.6209, 209.0858 59.7264, 250.83 66.83069999999999, 208.0173 58.7985, 160.9647 50.8049, 159.0115000000001 50.6209))" ;
		:geospatial_bounds_crs = "EPSG:4326" ;
		:geospatial_vertical_units = "m" ;
		:time_coverage_start = "2019-11-29T15:05:02Z" ;
		:time_coverage_end = "2020-04-27T08:29:22Z" ;
		:time_coverage_duration = "P149DT17H24M20S" ;
		:time_coverage_resolution = "P0DT0H42M21S" ;
		:date_issued = "2020-04-27T16:04:41Z" ;
		:date_modified = "2020-04-27T16:04:41Z" ;
		:argos_program_number = "11691" ;
		:creator_email = "michael.rehberg@alaska.gov" ;
		:first_uplink_date = "1575510820" ;
		:id = "5deb0b1d6321be14905284b8" ;
		:last_uplink_date = "1587997825" ;
		:ptt = "180473" ;
		:last_location_lat = "59.1356" ;
		:last_location_lon = "-151.4463" ;
		:last_location_date = "1587997825" ;
		:Conventions = "CF-1.6, ACDD-1.3" ;
		:acknowledgement = "NOAA IOOS, Axiom Data Science, Navy ONR,N OAA NMFS, Wildlife Computers, Argos" ;
		:creator_name = "Michael Rehberg" ;
		:creator_url = "https://www.adfg.alaska.gov/index.cfm?adfg=marinemammalprogram.stellerprogram" ;
		:infoUrl = "https://dev.axiomdatascience.com/?portal_id=99#search?type_group=all&query=habitat%20use%20of%20adult%20female%20steller&page=1" ;
		:institution = "Alaska Department of Fish and Game" ;
		:keywords = "atn,ioos,trajectory, steller sea lion" ;
		:license = "This animal telemery deployment data from Argos program 11691 and ptt 180473 is made available under the Open Database License: http://opendatacommons.org/licenses/odbl/1.0/. Any rights in individual contents of the database are licensed under the Database Contents License: http://opendatacommons.org/licenses/dbcl/1.0/" ;
		:metadata_link = "https://www.somelinkwhenwehaveacollectionpageat.NCEI.gov" ;
		:processing_level = "ATN DAC level 1 data prodcut [data levels yet to be explicitly documented[" ;
		:project = "Habitat Use of Adult Female Steller Sea Lions in the Endangered Western Distinct Population Segment, 2019-2020" ;
		:geospatial_lat_min = "50.6209" ;
		:geospatial_lat_max = "66.8307" ;
		:geospatial_lon_min = "-154.258" ;
		:geospatial_lon_max = "160.9647" ;
		:geospatial_vertical_min = "0.0" ;
		:geospatial_vertical_max = "0.0" ;
		:creator_country = "USA" ;
		:creator_institution = "Alaska Department of Fish and Game" ;
		:creator_sector = "gov_state" ;
		:date_metadata_modified = "2020-12-02T01:01:41Z" ;
		:instrument = "satellite telemetry tag" ;
		:platform = "animal" ;
		:platform_id = "5deb0b1d6321be14905284b8" ;
		:platform_name = "5deb0b1d6321be14905284b8" ;
		:platform_vocabulary = "https://mmisw.org/ont/ioos/platform" ;
		:program = "IOOS Animal Telemetry Network" ;
		:publisher_country = "USA" ;
		:publisher_institution = "US ATN DAC" ;
		:publisher_type = "institution" ;
		:vendor = "Wildlife Computers" ;
		:vendor_id = "5deb0b1d6321be14905284b8" ;
		:wmo_platform_code = "99nnnnn" ;
		:comment = "Flat Island, Alaska. Adult female with nursing pup (young-of-year). Brand X429. Mass not measured. \"SPLASH 10\" GPS location- and behavior-recording instrument glued to fur on top of the head." ;
		:sea_name = "North Pacific Ocean, Sea Okhotsk, and Bering Sea" ;
		:summary = "Wildlife Computers Splash 10 tag deployed on a Steller sea lion [Eumetopias jubatus] by Michael Rehberg in North Pacific Ocean, Sea Okhotsk, and Bering Sea from 2019-11-29 to 2020-04-27. PTT tag number 180473." ;
		:title = "Steller sea lion (Eumetopias jubatus) tag deployment from 2019-11-29 to 2020-04-27 in the North Pacific Ocean, Sea Okhotsk, and Bering Sea, ptt 180473" ;
		:history = "Mon Feb  8 14:31:10 2021: ncatted -a platform_groups,global,d,, Downloads/NCEI_test.2.nc Downloads/NCEI_test.3.nc\nMon Feb  8 14:28:47 2021: ncatted -a platform_category,global,d,, Downloads/NCEI_test.nc Downloads/NCEI_test.2.nc\nMon Feb  8 14:06:17 2021: ncks -x -v instrument,trajectory,deploy_id,type,comment,qartod_rollup_flag Downloads/atn_deployment_01.5.nc Downloads/atn_deployment_NCEI_test.nc\nnarrative description of ATN DAC processes for creating this file and sending to NCEI" ;
		:NCO = "4.7.2" ;
data:

 crs = _ ;

 ellipse_orientation = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, 74, 56, 57, 93, 50, 78, 67, 101, 113, _, _, _, _, _, _, _, 102, _, 
    _, 76, _, 167, _, _, 106, 106, 105, 88, _, 88, 88, _, 91, _, 92, 85, 125, 
    _, _, 101, _, _, 91, _, _, 89, _, 81, 84, 102, 88, 89, 89, 90, 91, 94, _, 
    _, _, 123, _, 97, _, 99, 90, 90, 89, 123, 116, 88, 90, 112, 91, 99, 96, 
    96, 82, 89, 84, 85, 85, 25, 41, 114, 72, 88, 87, 95, 92, 92, 87, 85, 85, 
    78, _, 81, 120, 65, 87, 88, 89, 113, 79, 166, 88, _, 106, 83, 104, 49, 
    47, _, _, _, _, _, _, _, _, _, _, _, 113, 91, 99, 100, _, 93, 78, 113, 
    84, 91, 112, _, 98, 94, 90, 96, 91, 51, 69, 72, 107, 87, 89, 86, 85, 84, 
    88, _, _, _, _, _, _, _, _, _, _, 72, _, _, _, 88, 86, 83, 84, 85, 86, 
    86, 89, 64, 84, 91, 90, 98, 95, 1, 58, 90, _, _, 90, _, _, _, 104, 90, 
    53, 73, 19, 58, 83, 171, 17, 70, 82, 89, 72, 106, 66, 50, _, 5, 102, 90, 
    79, 86, 80, 87, 87, _, _, _, _, _, _, _, _, _, _, 86, 153, 94, _, _, 80, 
    _, 96, 92, 110, 46, _, 97, 103, _, 44, _, 123, _, 86, 97, 88, 74, 89, 80, 
    75, 118, 126, 80, 96, _, _, 91, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, 61, _, 75, 80, 78, 61, 111, _, 90, 76, 84, 79, 81, 
    111, 91, 79, 82, 96, 113, 99, 89, _, 69, 71, _, _, _, _, _, _, _, _, _, 
    _, 29, 76, 48, 87, 76, 94, 90, 77, 120, 93, 70, 104, 70, 70, 98, 76, 86, 
    87, 139, 88, 100, 89, 106, 113, 53, 52, 84, 117, 81, 87, 83, 153, 153, 
    152, 85, 86, _, 98, _, _, 71, 77, 97, _, 75, _, 96, 133, 19, 94, 81, 139, 
    _, 83, _, 90, _, 98, _, 101, 94, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, 85, 85, _, _, _, 85, 148, _, _, _, _, 102, _, 105, 103, _, 68, 
    77, _, 161, 93, _, 87, 87, 94, 94, 98, 101, _, 79, 80, 76, _, 80, 80, 82, 
    _, _, _, _, _, _, _, 61, _, 158, _, 89, 94, 69, 121, 95, 93, 92, 92, 102, 
    93, _, _, _, _, 61, _, _, 58, _, 51, _, 87, _, 100, 86, 85, 89, 71, 72, 
    _, 72, 86, 110, 80, 84, 66, 86, 78, 98, 89, _, _, 86, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 85, 87, _, 88, _, 
    89, _, 92, 84, _, 89, 87, 99, 82, 85, 87, 92, _, _, _, 84, 38, _, _, 93, 
    _, 87, _, 114, 95, 114, 116, _, _, _, _, _, _, _, _, _, _, _, _, 49, 56, 
    87, 87, _, 83, 75, _, 107, 94, 74, 85, 137, 90, 82, 96, 83, _, _, 87, 
    124, 147, 94, 84, 109, 72, 101, 101, _, 69, 125, 92, 1, 91, 99, 101, 100, 
    100, 119, 176, 92, 87, 91, 92, 88, 88, _, _, _, 92, 92, _, 79, 79, 80, 
    93, 148, 106, 78, _, 81, 98, 100, 66, 79, 81, 79, 117, 79, 91, 91, _, 85, 
    88, 89, _, _, _, _, _, _, _, _, 17, _, _, _, _, _, 80, _, _, _, 119, _, 
    113, 105, _, _, _, 93, 100, 100, 70, _, 119, 89, _, 89, 113, _, 93, _, 
    89, 74, _, _, _, _, 77, 95, _, 91, _, 85, _, _, _, _, 106, _, 94, _, _, 
    _, _, 102, 78, 91, 90, 47, 106, 105, 78, 28, 105, 90, 140, 73, 98, 74, 
    75, 115, 80, 97, 96, 94, 87, 89, 117, _, _, _, _, _, _, _, _, _, _, 92, 
    22, 74, _, _, 82, _, 30, 76, 97, 45, 90, 68, 87, 69, 71, 101, 89, 90, 84, 
    91, 95, 91, 89, 129, _, _, _, _, _, _, _, 98, 98, 69, 55, 124, 96, 67, 
    87, 74, 84, 93, 79, 75, 79, 100, _, 68, 125, _, _, _, _, 128, 126, _, 95, 
    _, 130, 120, 97, 93, 56, 68, 108, 91, 176, 110, 99, 90, 51, 99, 91, 87, 
    117, _, _, 75, _, _, 84, 66, 138, 99, 109, 76, 81, 103, 98, 96, 73, 79, 
    105, 89, 97, 134, 75, 91, _, _, _, _, 89, 89, 81, 83, 81, 84, 83, _, _, 
    72, 75, 74, _, 8, _, _, 96, 84, 93, 75, _, 78, 74, _, 79, 85, _, 98, 76, 
    121, 73, 87, 89, 90, 94, _, _, 91, 99, 98, 90, 90, 86, _, 87, 4, 56, 85, 
    87, 88, 87, 107, 71, 89, 157, 1, 91, 91, _, _, 92, _, _, _, _, _, _, _, 
    84, _, 13, 106, 94, _, 90, 91, 89, 77, 111, 80, 73, _, 85, 95, 105, 59, 
    100, 79, 79, 111, 71, 78, 85, 95, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, 46, 80, 82, 56, 89, 160, 87, 88, 82, 67, 63, 99, 90, 90, 80, 85, 83, 
    112, 102, 130, 82, 80, 79, 82, 85, 86, 86, _, _, _, _, _, _, _, _, 82, 
    132, _, _, _, _, 102, 105, 90, 90, 106, 104, 96, 99, 97, 96, 94, 100, 90, 
    _, 86, _, 83, _, _, 79, 69, 72, 72, _, 76, _, 107, 104, 88, 100, 83, 113, 
    76, 111, 80, 103, 84, 79, 79, 112, 91, 89, _, 85, 175, _, _, 106, 91, 99, 
    82, 88, 89, 88, 80, 120, 12, 89, 3, 108, 177, 101, 76, 78, 85, _, 96, _, 
    80, _, 90, _, 102, _, 94, 105, _, _, _, _, _, 81, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 104, _, 88, _, _, 89, 
    89, 90, _, _, 86, 111, 96, 106, _, 103, 98, _, _, 81, 98, _, _, 69, _, 
    74, _, 106, 75, _, 109, _, 75, _, 93, _, 79, _, 83, 83, 110, 93, 93, _, 
    _, _, _, _, _, _, 93, 95, 99, 54, 78, 49, 132, 90, 104, 3, 99, 82, _, 86, 
    85, 89, 99, 73, 87, 89, 121, _, 125, _, 115, 90, 96, 92, 85, _, _, 84, _, 
    _, 85, 84, 26, 81, 86, _, 81, 84, _, 110, 100, _, 106, _, 99, _, _, _, _, 
    87, _, _, _, _, 56, 48, 71, 88, 42, 79, 78, 94, 90, 56, 65, 93, 87, 80, 
    113, _, 90, _, _, 94, _, 89, _, _, _, _, _, 90, 93, 92, _, _, _, _, _, _, 
    87, 84, 80, _, 88, _, 130, _, _, _, 86, 93, 112, 85, 83, 74, 83, 79, 99, 
    78, _, 77, 83, 67, 80, 91, 62, _, _, 83, _, _, _, 48, _, _, 81, 67, 79, 
    46, 122, 96, 83, 60, 88, 100, 73, 70, 88, 82, 114, 93, 92, 96, 87, 101, 
    74, 124, 79, _, 80, 4, _, 88, 9, 101, 95, 90, _, 92, _, _, 91, 90, 88, 
    92, _, _, _, _, _, 88, 48, _, _, _, _, 77, _, _, 79, _, _, _, 92, 93, _, 
    85, _, 89, 105, 75, 96, 103, 79, 78, _, 88, 102, _, _, 76, _, 79, _, 82, 
    _, _, _, _, _, 88, _, 66, _, _, 81, 86, _, _, 112, 134, 79, 101, 94, 114, 
    62, 57, 92, 129, 97, 76, 77, 83, 82, 116, 134, 126, 152, 109, 87, _, 78, 
    77, 98, 95, 82, 98, 76, 79, 79, 74, 95, 93, _, 161, 119, 97, 101, 98, 94, 
    88, 95, 112, 92, _, 81, 69, 82, _, _, _, 31, 33, _, 93, 144, 105, 80, 
    142, 115, 97, 73, 81, _, _, 87, 96, _, 78, 84, 88, _, _, 87, 74, 68, _, 
    89, 102, 101, _, 99, _, 96, 98, 93, 103, 102, 92, 92, 85, 95, 68, 25, 88, 
    _, 148, 145, 143, 75, 116, 91, 62, 67, 75, 118, 87, 80, 86, 81, 82, 176, 
    136, 104, _, _, _, _, _, _, 134, _, _, _, _, 75, 75, 96, 91, 92, 88, 83, 
    _, _, 91, 40, 88, 80, 87, 72, 65, 87, 159, 127, _, _, _, 136, _, _, _, _, 
    _, _, _, _, _, _, _, _, 58, 73, _, 86, 86, 66, 92, 167, 59, 87, 66, 96, 
    89, 78, 86, 122, 87, 81, 94, 111, 66, _, _, 75, 78, 68, 68, 80, 105, 79, 
    88, 77, 77, 95, 85, 95, 80, 75, 79, 75, 88, _, _, _, _, _, _, 97, _, 92, 
    91, 97, _, _, _, _, _, _, _, _, _, _, _, _, _, 79, 83, 89, 91, _, 100, 
    80, 87, 87, 85, 82, 81, _, 100, 151, _, 119, _, 92, 79, _, 79, 173, _, _, 
    69, 79, _, 51, 89, 91, _, _, _, 90, 87, 89, 91, 41, _, 110, 81, _, 105, 
    102, 100, _, _, _, 62, 88, 86, 77, 81, 92, 134, 74, 73, 10, 95, 20, 100, 
    93, 73, 72, 81, 76, 140, 92, 89, 106, 87, _, 96, _, _, _, _, 77, _, _, 
    68, _, 83, 85, 85, 85, 63, 63, 122, 85, _, 88, 120, 110, 76, 82, 101, _, 
    _, 19, 79, _, 102, _, _, 93, 118, 102, 50, 74, 86, _, _, _, _, _, 77, 76, 
    88, 108, 81, 114, 94, 114, 87, 80, 71, 89, 116, 105, 77, 83, 82, _, 87, 
    78, 97, 89, 123, 102, 108, _, _, _, _, _, _, _, _, _, _, 103, 101, 124, 
    _, 101, _, 134, 114, 103, 98, 176, 94, 99, _, 105, 100, 97, 93, 93, 103, 
    81, 76, _, 92, 84, 87, 94, 74, 80, _, _, _, 124, _, 21, 97, 72, 84, 91, 
    90, 90, 88, _, 93, _, _, _, _, 91, 98, 88, _, _, _, _, _, 91, 86, _, 89, 
    _, 78, 70, 5, _, 90, 175, 135, 92, 122, 67, 89, 158, _, 90, 90, 88, 87, 
    89, 89, 96, 94, _, 99, 2, 73, _, 79, 139, 83, 104, 123, 79, 89, 80, 100, 
    92, 81, 103, 98, 86, 84, 82, 81, 88, 82, _, _, 91, 110, 39, 79, _, 89, 
    62, 63, 99, 78, 94, 89, 72, 108, 88, 90, 84, 81, 79, 97, 79, 115, 107, 
    83, _, _, _, 90, _, 93, 78, 77, 99, _, 97, 95, 14, 104, _, _, 92, 74, _, 
    162, 79, 92, 100, 100, 64, _, 88, _, 79, _, 60, _, 78, 81, 83, 88, 90, _, 
    _, _, _, _, _, 17, _, 134, _, 147, 66, _, _, 118, _, 102, 126, 76, 34, _, 
    93, 90, 79, 100, 99, 59, _, 62, _, _, 149, 90, 114, 96, 108, 80, 90, 154, 
    102, 81, 82, 96, 137, _, _, _, _, _, _, _, _, _, _, _, 79, 128, _, 80, 
    82, _, 96, 97, 77, _, _, _, _, _, _, _, _, _, _, 51, _, _, 74, _, 107, 
    102, _, 93, _, 85, _, 86, 86, 120, _, 84, _, 86, _, 87, _, _, 71, 89, 85, 
    86, 95, 80, 84, 88, _, 123, _, _, 162, 67, 93, 83, 89, _, 32, _, 59, 175, 
    89, 87, 89, 90, 31, 79, 96, 86, 116, 95, 41, 80, 108, 116, _, _, 93, 48, 
    89, 80, 68, 20, 86, 118, _, 91, 90, _, 104, 96, 90, 30, 86, 87, 72, 103, 
    83, _, 79, 93, _, 89, 88, 89, _, 85, 79, _, _, _, _, 8, _, 77, _, 89, _, 
    106, 94, 91, 5, 87, _, 103, 91, 96, 85, 87, 109, 76, 77, 82, 92, 93, 91, 
    85, 87, 89, _, _, _, _, _, 127, _, 92, 62, 81, 85, _, _, _, _, _, _, _, 
    71, 87, 101, 77, 55, 84, 132, 56, _, 57, 92, 80, 122, 90, 103, 80, 89, 
    89, 93, _, _, 89, 92, 112, _, _, _, _, _, 121, 91, 97, 89, _, 89, 88, 96, 
    77, 89, 119, 94, 50, 73, 105, 66, 87, _, _, 66, 82, 89, 88, 126, 76, 121, 
    117, 114, _, _, _, _, _, _, 79, 82, 88, 103, 91, 100, 93, 89, 173, 79, 
    81, 78, 71, 71, _, 83, _, 85, _, 116, _, _, _, _, _, _, _, _, 90, 30, 74, 
    80, _, _, _, 66, 154, 77, 77, 74, 66, _, _, _, _, 80, 79, 60, _, 75, 90, 
    107, _, _, 110, 30, 89, 88, _, 104, 91, 89, _, 101, 96, _, _, 93, 98, 88, 
    88, 102, _, _, _, _, 101, 93, _, 78, 81, 83, 85, 85, _, 89, 90, 89, 137, 
    121, 104, 96, 74, 81, 66, 80, 85, 77, 98, _, 118, 126, _, _, _, 86, _, _, 
    _, 86, _, 82, _, 149, _, _, _, _, 55, 56, _, 143, _, 107, _, _, 72, _, 
    104, 43, _, 158, 91, _, 91, 89, 85, 138, _, _, 71, _, 73, 88, 94, 92, 71, 
    91, 92, 77, 129, 90, 90, 100, _, 88, _, 95, 68, 87, _, _, 89, 115, _, 96, 
    96, _, _, _, 94, 94, 93, 100, 88, _, _, _, _, _, _, 93, 95, 92, 80, 111, 
    103, 72, 105, 69, 84, 86, 103, 104, 81, 98, 84, 104, _, 66, 86, 87, 120, 
    85, 90, 87, 127, _, _, _, 75, 73, 88, 61, 95, 90, 92, _, _, 50, 88, 116, 
    110, 91, 68, 88, 105, 81, 87, 86, 87, 113, _, _, 80, 114, _, 92, 98, _, 
    101, 99, _, 123, 58, 73, 103, 105, 71, 92, 94, _, 90, _, _, _, 97, 97, 
    93, 90, 62, 68, _, 77, 83, 160, 64, 78, 136, 101, _, 96, 106, 93, _, 90, 
    71, 78, 89, _, 82, 91, 74, _, 84, 89, 90, 101, _, _, _, _, 88, 70, _, _, 
    _, 67, _, _, 69, 91, 104, 102, _, _, _, 58, _, _, 109, _, 101, 92, _, 85, 
    _, _, 62, _, _, 90, 98, _, 114, 95, _, 92, 85, _, 93, 77, 78, 80, 83, _, 
    83, _, 69, 81, _, 116, 106, 100, 89, 77, 54, 100, 80, 79, 93, 88, _, 98, 
    99, _, 66, 86, 99, _, 95, _, 138, _, _, _, _, _, _, _, 92, 84, 92, _, _, 
    _, _, 69, 115, 107, 94, 81, _, 66, _, 98, 97, 56, 76, 77, 61, 101, 60, 
    79, 87, 87, 92, 118, 84, 107, 117, 91, _, _, _, _, _, _, _, 77, 80, 77, 
    101, 73, 81, 55, _, 96, 61, _, _, 79, 91, 89, _, 110, 83, 87, 106, 90, _, 
    _, _, _, _, _, _, _, _, _, _, _, 70, _, _, 75, 81, 85, 83, 86, 83, 85, 
    87, 92, 0, 90, 168, 82, 78, 82, 84, 83, 171, 58, 105, 91, 88, 33, 67, 71, 
    81, 178, 153, 73, 77, 94, 80, 44, 53, 87, 88, 89, 115, 104, 75, 74, 67, 
    82, 106, 97, 93, 116, 87, _, _, _, _, _, _, _, _, _, _, 34, 73, 14, 71, 
    90, 89, 3, _, 88, 80, 88, 90, 94, 99, 67, 88, 137, 79, 70, 80, _, 96, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, 77, 123, _, _, 106, _, _, 93, 85, 85, 
    66, 97, 93, 71, 104, 80, 96, 90, 86, 56, 83, 49, 103, 108, 75, 81, 77, 
    98, 52, _, 67, 84, _, _, _, _, _, _, 94, _, 99, _, 101, 97, 79, 63, _, 
    68, 116, _, 96, 95, _, 111, _, 77, _, 82, _, 86, 79, 81, _, 89, 90, 87, 
    87, 90, 90, _, _, _, _, _, 93, _, _, 93, 90, _, _, 94, 103, 124, 114, 76, 
    96, 107, 109, 179, 90, 90, 90, 102, _, _, _, _, _, _, _, 43, 51, _, _, 
    85, 70, 70, 22, 74, 67, _, 118, 106, 99, 87, 80, _, 83, _, 84, _, _, 22, 
    82, _, 89, 58, _, _, _, _, 84, 105, 173, 80, 172, 89, 64, 22, 109, 91, 
    100, 86, 72, 74, 103, 80, 88, 82, 96, 93, 95, 93, 98, 76, 89, _, _, _, 
    79, _, 87, _, 87, 34, 65, 67, 90, 80, 83, _, 84, 99, 112, 70, 83, 78, _, 
    80, 103, 79, 83, 169, 117, 109, 31, _, _, _, _, _, _, _, _, _, _, 139, 
    57, _, 42, 71, 37, 88, _, 77, 108, _, 91, 51, 100, 84, 109, 83, 78, 86, 
    _, 78, 81, _, 81, 88, _, _, _, _, _, _, _, _, _, 103, 87, 91, 88, _, 75, 
    _, 82, _, 108, 124, 103, _, 73, 78, 80, _, 45, 98, 61, 79, 87, 78, 106, 
    83, _, 80, _, 59, 67, 89, 90, 89, _, 86, _, _, _, _, _, 178, _, 75, _, _, 
    _, _, _, _, _, _, _, 64, 122, 78, 89, 101, 93, _, 93, _, _, 68, 63, 179, 
    90, _, _, 53, 62, _, 95, 78, _, _, 76, _, 87, 88, 74, 78, 123, 114, 101, 
    _, _, 173, 172, 1, 89, 91, 40, 27, 94, 140, _, 90, _, _, 89, 79, 100, 97, 
    73, 41, 80, 98, 91, 68, 87, 90, 41, 15, 90, _, 86, _, 119, 105, _, _, _, 
    96, 89, 88, 88, 111, 110, 76, 122, 91, 95, 96, 90, 85, 85, 40, 101, 100, 
    100, 100, _, 95, 95, 115, 96, 90, _, _, _, _, _, _, _, _, 66, 66, _, 68, 
    _, _, _, 93, 93, 92, 92, _, 87, 83, 122, 76, 8, 87, 86, 66, 86, 46, 87, 
    90, 90, _, _, 90, 114, 93, 85, _, 91, 83, _, _, 82, 80, 93, 96, 90, 93, 
    86, 89, 90, 100, _, 81, 61, 76, 88, 62, 85, 62, 101, 72, 81, 92, 78, 90, 
    89, 109, 42, 60, _, _, _, _, _, _, 72, 85, 85, _, _, 72, 79, _, _, 79, 
    132, 115, 99, _, 99, _, _, 62, _, 78, 71, _, 49, 65, _, 103, _, 81, 75, 
    _, _, _, _, _, _, _, _, _, 92, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, 82, 84, _, _, 77, _, 88, _, 74, 100, 90, 85, 88, 88, 87, 86, 79, 75, 
    115, 83, 88, _, 91, 64, 101, 70, 131, _, 76, _, _, 66, _, 82, 42, 99, 
    123, 68, 78, 103, 62, 80, 75, _, 73, 88, 98, 143, _, _, 153, 125, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, 68, _, _, 49, 88, 95, 92, 91, 90, 
    94, 94, 88, 88, 69, 82, 74, 89, 86, 76, 100, 120, _, 89, _, _, _, _, 89, 
    89, 101, 95, 92, 102, 72, 169, _, 110, 86, 87, 101, _, _, 94, 89, 79, _, 
    92, _, _, 89, 91, 89, 89, 130, 97, 77, _, 65, _, _, 99, 72, _, _, 115, _, 
    65, 86, 32, 95, 87, 69, 81, 43, 143, 109, 72, 93, 104, 89, 90, 107, _, 
    111, 90, 89, _, 91, 92, 100, 110, 96, 94, 90, 93, 94, 94, _, _, 93, _, 
    93, 93, _, 93, 92, 60, _, 82, _, 84, 88, 89, 17, 88, 111, 102, 91, 69, 
    98, 97, 95, 73, 85, 84, 64, 99, 93, 92, 126, 58, 56, 80, 79, 91, 120, 91, 
    _, _, 100, 72, 6, 131, 92, 92, _, _, _, 93, 79, 86, 93, 101, 84, 96, 94, 
    89, 88, 83, 79, 79, 91, 129, 95, 91, _, 139, 91, 92, 167, 71, 112, 109, 
    79, 90, 92, 91, _, 73, _, _, _, 87, 75, 75, 79, _, 78, _, 79, _, 101, 77, 
    70, _, 131, 95, 91, 102, 93, 69, 71, 131, 70, _, _, _, 96, _, _, 90, _, 
    _, _, _, 91, 79, 79, 72, _, 75, 58, 81, 82, 143, _, _, 93, 80, 80, 79, 
    89, 108, 100, 48, _, 77, 67, 109, 97, 129, 93, 85, 86, 96, 101, 32, 89, 
    89, 89, 89, 94, 63, 76, 90, 98, _, _, _, _, 133, 128, 36, 88, 91, 84, _, 
    _, _, _, 90, 93, 93, 139, 75, 49, 86, 81, 110, 101, 108, _, 79, 84, 104, 
    101, 95, 78, 94, 84, 77, _, 150, 86, 104, _, 149, _, 121, 119, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, 81, _, _, _, 73, _, 86, _, 92, 91, _, 124, 
    77, 110, 76, 89, 110, 103, 77, 89, 52, 144, 63, 82, 152, 80, 97, 87, 115, 
    85, 49, _, _, _, _, 113, _, 56, _, 89, 75, 73, 74, 104, 82, 107, 70, 80, 
    77, 79, 88, 110, 79, 84, 85, 91, 89, 49, 75, 94, _, _, _, _, _, _, _, _, 
    57, _, 88, _, 88, 88, _, _, 88, 87, 98, _, _, 100, 77, _, 78, _, 103, 85, 
    78, _, 96, _, 99, 94, 109, 93, 91, _, 15, _, 27, _, _, 130, 89, 87, _, _, 
    102, _, _, 106, 63, _, 77, _, _, 84, 84, _, _, 100, 90, 97, _, 100, _, _, 
    99, 91, 88, 73, 77, _, _, _, 116, 158, _, 77, 84, _, 72, 87, 114, 99, _, 
    93, _, _, _, 74, 86, _, 88, 78, 86, 89, _, 59, 68, _, _, _, 86, 20, _, _, 
    86, _, _, 93, _, 123, _, 81, _, 100, 66, 86, 96, 87, 101, 118, 161, 107, 
    96, 82, 118, _, _, _, _, 88, 88, _, 92, 93, 109, _, 92, _, 86, _, 86, 99, 
    114, 79, 72, 71, 98, 81, 83, 98, _, 90, 90, _, _, _, 160, _, _, 102, 45, 
    89, 110, 174, _, _, _, _, _, _, 152, _, 143, 140, 124, _, _, 78, 78, 78, 
    103, 99, 99, 96, 69, 85, _, 76, _, 77, _, _, 81, _, _, 72, 72, 75, 65, _, 
    83, 86, 98, 91, 96, 107, _, 101, 106, _, _, _, _, _, 80, _, 8, _, 91, 80, 
    75, 68, 78, 102, 102, 121, 113, 80, _, 89, 86, _, 82, 89, 85, 84, 82, 92, 
    87, 159, 93, 93, 134, 83, 88, 117, 89, 151, 90, 86, 100, 115, 60, 45, 78, 
    _, 82, 83, 108, 100, 87, 87, 96, _, _, _, _, 93, _, _, 86, 91, 98, 77, 
    77, 83, 44, 20, _, _, _, _, 93, 74, _, 102, 102, 6, 69, 94, 21, 71, 86, 
    89, 45, 55, 92, 92, 84, 113, 105, 60, 63, 81, 107, 126, 78, 81, 81, 111, 
    110, 156, 73, 79, _, 70, 85, 85, 101, 115, _, 90, 89, 89, 113, 106, 98, 
    102, 102, 101, 75, 82, 118, 93, 90, 93, _, 91, 22, _, 176, 98, _, _, 77, 
    79, 85, 75, 86, 113, 106, 85, _, 88, 91, 78, 79, 87, 88, 99, 122, 95, _, 
    137, _, _, _, 88, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 66, 47, _, 
    81, 98, 8, 86, 121, 131, 76, 57, 90, 118, _, 105, 75, _, _, 69, _, 81, _, 
    111, 91, _, 90, 83, 88, 96, _, _, 107, _, 25, _, _, _, _, 52, 107, 106, 
    104, 33, 63, 91, _, 152, _, 72, _, 81, 13, 100, 71, 42, _, 139, 71, 83, 
    90, 55, 55, _, _, 79, 95, 90, 82, 92, 90, 89, 101, 133, 88, 19, 61, 150, 
    74, 87, 73, 81, 41, 89, 92, 59, 77, 54, 43, 101, 89, 79, 98, 81, 87, 50, 
    103, 92, 164, 81, 69, _, 83, 80, 89, 77, _, 69, 72, _, _, _, _, 84, _, _, 
    90, _, _, 151, _, _, 96, _, 86, _, _, _, _, _, 89, 85, _, 96, _, _, _, 
    86, 85, 39, 106, 124, _, 142, 119, 93, 93, 92, 74, _, _, 66, _, _, _, _, 
    75, 81, _, 86, 87, _, 105, 91, _, 102, 101, 100, 35, 78, 80, 83, 85, 83, 
    85, _, _, 90, 95, _, _, 81, 86, 104, 99, 99, 81, 89, 135, 158, 97, _, _, 
    _, 103, 57, 84, 87, 87, 92, 92, 91, 54, 70, 86, 86, 68, 86, 80, 81, 125, 
    110, 106, 101, 85, 103, 82, 83, 56, _, _, 83, 87, _, _, 83, 129, 115, 79, 
    99, _, 88, 83, _, 95, _, _, _, 70, 67, 88, 108, 118, 104, 169, 89, 108, 
    87, 111, 112, 127, 10, 98, 79, 91, 82, 81, _, 85, _, 89, 103, _, _, _, 
    68, _, 66, _, _, 103, 98, 99, _, 9, _, 14, _, _, _, _, _, _, _, 37, _, 
    132, _, 66, 68, 76, 84, 83, 77, 88, 83, 114, 65, 82, 85, 104, 80, 82, 80, 
    _, 86, 150, 137, 103, _, 97, 49, _, 177, 88, 88, 99, _, _, _, _, _, _, _, 
    _, _, _, 126, 47, 55, 29, 79, 81, 59, 66, 81, 51, 105, 151, 69, 87, 89, 
    103, 76, 78, 73, 85, 98, 99, 109, 76, 67, _, _, 79, 85, 148, _, 97, 95, 
    71, _, 85, _, _, _, 91, 155, _, _, 86, 73, _, 98, 90, _, 89, 160, 120, 
    86, 90, 101, 51, 90, 90, 99, 107, 93, 94, 99, 89, 76, 86, 125, _, 103, 
    118, 125, 104, 80, 88, 86, _, 74, 89, 73, 120, 61, 79, 88, 88, _, 88, 90, 
    35, _, _, 82, _, _, _, _, _, _, _, _, 73, 42, 77, 88, _, _, 75, 85, 89, 
    87, 155, 68, 94, 100, 94, 90, 10, _, 57, 85, 38, _, _, 68, _, _, 84, 83, 
    63, 85, 34, 90, 90, _, _, _, _, _, _, _, _, 91, _, _, _, 79, 154, 74, 
    146, 149, 62, 75, 57, 77, 88, 98, 91, 86, 123, 89, 78, 75, 135, 78, 88, 
    _, 104, 113, 102, 89, _, 88, _, 40, 87, 82, 88, 96, 94, 100, 97, 95, _, 
    97, _, 91, 63, 90, 151, 107, 109, 72, 76, 89, 88, 89, 99, 90, 75, 99, 79, 
    111, 88, 98, 82, 104, 90, 90, 76, 87, 80, 91, 86, 15, _, 21, 55, 114, _, 
    _, _, _, _, _, _, 112, 69, 86, _, 89, 89, 62, 78, 85, 84, 91, 91, 80, 89, 
    98, 96, 93, 88, 81, 82, 93, 104, 103, 93, 92, 109, 92, 90, 100, 122, 112, 
    107, 80, 83, _, _, 79, 81, 80, 110, 97, 90, 147, 106, 96, 115, 101, 84, 
    53, 70, 76, 80, 82, 87, _, 89, 126, 13, 89, 72, _, _, _, _, 72, _, _, _, 
    171, 75, 105, _, 117, 84, 100, 110, 95, 90, 87, _, 87, 141, 123, _, 93, 
    85, 88, 75, 33, 64, 125, 95, 67, 89, 101, 68, 6, 97, 97, _, _, 100, 78, 
    80, 83, 81, _, 93, 92, 96, 88, 92, _, _, _, _, _, 81, _, _, 75, 84, 138, 
    93, 80, _, _, _, 116, 124, 114, _, _, 95, 110, 167, 93, 90, 100, 147, 98, 
    117, 105, 99, 98, 96, 75, 111, _, 88, _, 88, _, 86, 72, 86, 119, 94, _, 
    _, 109, _, _, _, _, _, _, 125, 95, 136, 58, 86, 99, 100, 100, 60, 92, 54, 
    _, _, 99, 84, 90, 89, 66, 71, 79, _, 81, 154, 113, 82, _, _, _, _, 52, 
    107, _, 79, 90, _, 92, _, _, _, _, 74, 77, _, _, 83, _, 97, _, _, 96, 
    177, 86, _, 87, _, 101, 97, _, 87, 91, 93, 88, 88, 51, 158, 78, 85, 87, 
    _, 106, 84, 87, _, 26, 75, 82, 88, 101, 28, 98, 91, 90, _, 91, 66, 118, 
    96, 77, 79, _, 72, 80, 93, 68, 85, _, _, 88, _, _, 115, 73, 161, 70, _, 
    _, _, _, 69, _, _, 88, 53, 60, 61, 103, 99, 93, 117, _, 90, 78, 97, 94, 
    80, 78, 97, _, 92, _, 105, 95, 93, 101, 101, _, 85, 41, 78, _, 94, 89, 
    109, 106, 121, _, _, 109, 128, 99, 97, 92, 142, 94, 85, 102, 52, 64, _, 
    75, 75, 77, 83, 87, 44, 102, 85, _, 27, _, _, _, 76, 68, 96, 98, 95, 164, 
    106, 141, 138, 44, _, 77, 84, _, 72, _, _, _, 86, _, 107, _, 97, 90, 90, 
    72, 91, _, _, _, _, _, _, _, 80, 92, _, _, 88, 90, 99, 73, 108, 120, 90, 
    90, 68, 82, 81, 58, 78, 70, 76, 74, 99, 90, 94, 96, 89, 89, _, _, _, _, 
    120, 120, 99, 97, 119, 96, _, 178, _, 91, 93, _, 156, 122, 61, 123, 103, 
    _, 92, _, _, _, _, _, _, _, 23, _, _, 54, 79, _, 62, 92, 86, 46, 90, 100, 
    100, 74, 85, 92, 82, 90, 89, 118, 98, 98, _, _, _, _, _, _, 108, _, 83, 
    76, 68, 83, 105, 102, _, 95, 96, 123, 97, _, 84, 4, 4, _, 13, 79, 66, 83, 
    172, 96, 73, 52, 117, 118, 119, 99, 95, 83, 88, 89, 91, 86, 117, _, 121, 
    162, _, _, _, 120, _, 77, 78, 98, 58, 89, 79, 21, 85, _, 79, 88, 142, _, 
    106, _, 110, _, 67, _, _, 102, _, 91, _, 96, 99, _, 160, 84, 98, 89, 96, 
    111, 89, 98, 77, 81, 82, 89, 89, 91, 79, 85, 53, 43, 111, 92, 100, 85, 
    65, 82, 71, 11, 10, 44, 85, 76, 87, 86, 86, 57, 110, 119, 93, 89, 110, 
    63, 92, 81, 90, 83, 80, 76, 81, 77 ;

 error_radius = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    336, 272, 501, 412, 341, 512, 145, 164, 1681, _, _, _, _, _, _, _, 2039, 
    _, _, 1906, _, 1103, _, _, 1433, 1322, 1080, 544, _, 735, 1301, _, 1308, 
    _, 1394, 367, 923, _, _, 1523, _, _, 1858, _, _, 2780, _, 2790, 609, 379, 
    650, 1037, 1033, 861, 1003, 907, _, _, _, 1806, _, 2665, _, 2685, 1975, 
    1582, 2017, 1043, 1241, 362, 1448, 1410, 6513, 3578, 4272, 897, 896, 
    3268, 1197, 1306, 1344, 1023, 1142, 633, 227, 1052, 1146, 951, 1387, 
    1466, 960, 509, 520, 948, _, 1248, 813, 720, 377, 2013, 2130, 1327, 3149, 
    4271, 563, _, 466, 273, 244, 343, 1125, _, _, _, _, _, _, _, _, _, _, _, 
    270, 439, 1627, 1238, _, 1878, 300, 277, 277, 12332, 2024, _, 3207, 3648, 
    2487, 293, 1057, 205, 124, 314, 1936, 428, 297, 412, 175, 467, 5677, _, 
    _, _, _, _, _, _, _, _, _, 162, _, _, _, 1166, 938, 1338, 1567, 1602, 
    1735, 1787, 144, 1366, 1398, 1087, 455, 1234, 1525, 1565, 553, 699, _, _, 
    1509, _, _, _, 3550, 3449, 772, 1096, 411, 1698, 453, 1474, 1282, 357, 
    321, 2360, 152, 381, 316, 456, _, 970, 393, 1546, 1543, 2305, 4357, 4057, 
    2983, _, _, _, _, _, _, _, _, _, _, 5892, 381, 813, _, _, 1451, _, 2334, 
    580, 793, 189, _, 569, 259, _, 623, _, 1513, _, 227, 340, 1669, 179, 904, 
    1139, 174, 169, 657, 271, 431, _, _, 2751, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, 7992, _, 4953, 5405, 4667, 804, 413, _, 
    1227, 264, 834, 931, 461, 208, 869, 301, 583, 3779, 3957, 230, 1335, _, 
    1016, 937, _, _, _, _, _, _, _, _, _, _, 382, 169, 283, 1088, 210, 195, 
    908, 936, 564, 889, 148, 232, 241, 188, 223, 300, 341, 274, 1394, 161, 
    202, 702, 293, 735, 3533, 4072, 175, 238, 1180, 1224, 1164, 1422, 1442, 
    1439, 171, 260, _, 2590, _, _, 688, 478, 337, _, 324, _, 848, 564, 430, 
    1884, 261, 525, _, 556, _, 1274, _, 623, _, 440, 1123, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, 3650, 2181, _, _, _, 2430, 881, _, _, _, _, 
    1316, _, 1089, 264, _, 565, 497, _, 536, 126, _, 741, 718, 790, 954, 
    3469, 1534, _, 3892, 3146, 1160, _, 3918, 3138, 5464, _, _, _, _, _, _, 
    _, 8634, _, 931, _, 1207, 902, 174, 270, 497, 728, 707, 1043, 967, 215, 
    _, _, _, _, 3488, _, _, 450, _, 1684, _, 3622, _, 5206, 944, 622, 3312, 
    2403, 728, _, 1134, 751, 1062, 418, 1332, 1308, 489, 431, 187, 1502, _, 
    _, 1919, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, 267, 2052, _, 1529, _, 1076, _, 999, 305, _, 1711, 1280, 991, 
    389, 558, 878, 192, _, _, _, 810, 975, _, _, 770, _, 286, _, 346, 583, 
    1417, 1635, _, _, _, _, _, _, _, _, _, _, _, _, 5195, 2542, 421, 699, _, 
    776, 714, _, 503, 908, 243, 1190, 933, 1245, 756, 459, 179, _, _, 1284, 
    1237, 512, 1030, 215, 212, 727, 3747, 2967, _, 240, 834, 1016, 680, 2210, 
    1235, 812, 846, 867, 1010, 669, 700, 508, 4247, 4299, 4068, 4027, _, _, 
    _, 1648, 2095, _, 5229, 4173, 3457, 1040, 1221, 521, 762, _, 230, 206, 
    2020, 1077, 233, 1502, 805, 708, 735, 296, 607, _, 1693, 2010, 1036, _, 
    _, _, _, _, _, _, _, 800, _, _, _, _, _, 1738, _, _, _, 1137, _, 1131, 
    888, _, _, _, 1432, 1211, 1243, 308, _, 769, 1103, _, 1364, 1877, _, 
    5195, _, 5169, 336, _, _, _, _, 1088, 1801, _, 5793, _, 1427, _, _, _, _, 
    420, _, 1418, _, _, _, _, 1475, 685, 368, 3272, 600, 231, 183, 234, 391, 
    196, 236, 812, 514, 1345, 280, 361, 379, 580, 214, 457, 195, 867, 1993, 
    415, _, _, _, _, _, _, _, _, _, _, 3195, 3624, 886, _, _, 1500, _, 2287, 
    473, 193, 3567, 297, 222, 1482, 456, 164, 162, 1291, 158, 1590, 269, 145, 
    229, 1097, 1263, _, _, _, _, _, _, _, 4619, 3297, 7022, 3000, 745, 988, 
    637, 817, 278, 687, 512, 145, 312, 576, 404, _, 334, 547, _, _, _, _, 
    945, 999, _, 1721, _, 2058, 2997, 307, 2380, 1163, 782, 269, 758, 591, 
    145, 174, 1287, 294, 146, 3244, 3818, 1200, _, _, 810, _, _, 7614, 4839, 
    643, 684, 324, 260, 208, 490, 755, 779, 2767, 1001, 929, 1372, 282, 2446, 
    235, 1823, _, _, _, _, 1661, 6473, 5875, 922, 892, 1216, 1335, _, _, 
    1117, 1070, 1065, _, 1036, _, _, 1074, 1222, 755, 1318, _, 1199, 1269, _, 
    1200, 1693, _, 184, 775, 680, 206, 1550, 1689, 528, 659, _, _, 4982, 165, 
    446, 872, 638, 648, _, 383, 894, 619, 391, 440, 1509, 1667, 1128, 175, 
    837, 1853, 1417, 1485, 1404, _, _, 1623, _, _, _, _, _, _, 17948, 2900, 
    _, 1046, 460, 1642, _, 260, 517, 2235, 598, 725, 221, 329, _, 1141, 1288, 
    390, 378, 206, 559, 246, 772, 420, 1416, 1498, 3370, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, 299, 623, 749, 291, 1967, 961, 147, 377, 256, 250, 
    1243, 133, 245, 381, 293, 216, 468, 628, 728, 761, 1484, 1529, 4713, 
    4048, 3687, 2172, 2294, _, _, _, _, _, _, _, _, 428, 1065, _, _, _, _, 
    172, 148, 476, 478, 908, 1012, 916, 812, 1034, 1264, 1531, 159, 863, _, 
    1188, _, 1671, _, _, 2168, 943, 1070, 1080, _, 1307, _, 564, 465, 661, 
    666, 563, 410, 1921, 1256, 2137, 1253, 3367, 662, 1092, 217, 701, 1341, 
    _, 3399, 755, _, _, 772, 1939, 2337, 823, 2242, 5341, 1664, 533, 315, 
    191, 485, 208, 171, 1481, 751, 262, 306, 385, _, 975, _, 4421, _, 357, _, 
    146, _, 465, 968, _, _, _, _, _, 7218, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, 324, _, 2044, _, _, 181, 672, 
    788, _, _, 483, 566, 138, 295, _, 396, 223, _, _, 442, 178, _, _, 417, _, 
    523, _, 325, 245, _, 1040, _, 237, _, 208, _, 377, _, 685, 660, 1474, 
    1686, 1953, _, _, _, _, _, _, _, 4014, 3536, 3470, 1580, 799, 1400, 1801, 
    213, 1154, 248, 429, 1209, _, 2394, 434, 3480, 1621, 320, 140, 654, 593, 
    _, 857, _, 940, 884, 1090, 1257, 1469, _, _, 2609, _, _, 2780, 2865, 
    5158, 3239, 7429, _, 1677, 1059, _, 2087, 5257, _, 1656, _, 939, _, _, _, 
    _, 2153, _, _, _, _, 362, 3219, 747, 1022, 9444, 197, 1066, 167, 917, 
    243, 188, 462, 3561, 1170, 181, _, 880, _, _, 397, _, 2723, _, _, _, _, 
    _, 5145, 548, 875, _, _, _, _, _, _, 2043, 3348, 1305, _, 273, _, 428, _, 
    _, _, 142, 173, 246, 350, 147, 334, 352, 212, 158, 183, _, 1009, 230, 
    2307, 159, 183, 626, _, _, 2729, _, _, _, 2582, _, _, 541, 294, 259, 535, 
    730, 570, 238, 336, 1556, 355, 184, 154, 603, 726, 964, 258, 126, 584, 
    976, 674, 3594, 2608, 4954, _, 5922, 2584, _, 3079, 779, 256, 145, 992, 
    _, 1070, _, _, 1458, 1680, 1751, 1925, _, _, _, _, _, 2527, 537, _, _, _, 
    _, 3182, _, _, 4146, _, _, _, 247, 1136, _, 3095, _, 1592, 904, 750, 610, 
    844, 312, 563, _, 1065, 410, _, _, 1666, _, 1732, _, 972, _, _, _, _, _, 
    1619, _, 2574, _, _, 475, 925, _, _, 468, 383, 319, 547, 153, 623, 360, 
    671, 542, 2420, 1267, 1403, 868, 675, 834, 1291, 531, 667, 247, 735, 
    2127, _, 366, 731, 982, 646, 474, 598, 422, 487, 1950, 1755, 2312, 2281, 
    _, 2339, 375, 534, 541, 761, 1061, 1366, 266, 3055, 914, _, 13088, 16481, 
    12879, _, _, _, 1353, 1352, _, 238, 554, 745, 323, 592, 993, 1867, 355, 
    1772, _, _, 5842, 845, _, 389, 476, 1653, _, _, 2102, 2367, 828, _, 9294, 
    5530, 3001, _, 3183, _, 1764, 2353, 1799, 316, 185, 737, 1453, 3995, 
    4942, 550, 723, 1717, _, 1824, 841, 867, 576, 423, 214, 1638, 395, 764, 
    462, 649, 1002, 2762, 134, 324, 421, 1272, 796, _, _, _, _, _, _, 1389, 
    _, _, _, _, 2279, 3999, 1092, 835, 996, 957, 881, _, _, 687, 220, 689, 
    430, 165, 301, 201, 864, 1262, 2624, _, _, _, 1007, _, _, _, _, _, _, _, 
    _, _, _, _, _, 574, 1432, _, 3638, 152, 535, 315, 651, 1666, 3425, 884, 
    186, 580, 223, 551, 203, 201, 220, 641, 156, 609, _, _, 2047, 2429, 2248, 
    2234, 14804, 8890, 1678, 2429, 3437, 5503, 2466, 692, 287, 309, 613, 256, 
    775, 1378, _, _, _, _, _, _, 2584, _, 406, 3059, 1964, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, 2705, 226, 697, 623, _, 180, 1087, 1535, 2628, 4223, 
    1243, 1185, _, 1031, 630, _, 329, _, 934, 814, _, 839, 392, _, _, 471, 
    542, _, 299, 466, 1333, _, _, _, 3265, 2849, 2892, 2782, 1044, _, 716, 
    1133, _, 1047, 1049, 1158, _, _, _, 166, 392, 1119, 715, 907, 1076, 673, 
    208, 376, 972, 413, 199, 265, 144, 210, 200, 326, 1003, 450, 309, 514, 
    212, 1261, _, 8323, _, _, _, _, 1049, _, _, 3477, _, 363, 539, 730, 808, 
    705, 678, 820, 220, _, 626, 444, 688, 429, 821, 765, _, _, 368, 537, _, 
    1949, _, _, 4866, 1390, 1469, 347, 698, 1089, _, _, _, _, _, 5597, 401, 
    1746, 1401, 128, 429, 1409, 384, 375, 280, 260, 1822, 1343, 140, 172, 
    668, 3315, _, 4569, 414, 1608, 5961, 768, 2400, 2959, _, _, _, _, _, _, 
    _, _, _, _, 4608, 4141, 292, _, 587, _, 582, 794, 2212, 3262, 603, 767, 
    951, _, 695, 5004, 5907, 2425, 2502, 156, 1411, 426, _, 295, 609, 528, 
    249, 1049, 1725, _, _, _, 3114, _, 2589, 6063, 2369, 1857, 860, 1272, 
    1353, 1530, _, 1279, _, _, _, _, 2831, 3006, 2624, _, _, _, _, _, 421, 
    798, _, 2484, _, 168, 299, 368, _, 599, 690, 404, 211, 391, 301, 506, 
    203, _, 896, 695, 441, 566, 691, 2175, 1863, 1465, _, 184, 1824, 925, _, 
    1654, 686, 212, 353, 239, 169, 581, 694, 597, 378, 166, 498, 1753, 2056, 
    2767, 278, 233, 741, 712, _, _, 6379, 189, 1536, 159, _, 869, 381, 392, 
    919, 1580, 174, 447, 235, 706, 211, 319, 680, 1774, 385, 133, 2338, 1281, 
    1966, 511, _, _, _, 4021, _, 7167, 4503, 1977, 890, _, 1664, 1901, 912, 
    418, _, _, 1023, 1787, _, 1534, 2257, 2528, 1087, 1113, 591, _, 2205, _, 
    1401, _, 270, _, 801, 443, 270, 1048, 400, _, _, _, _, _, _, 1831, _, 
    1276, _, 1647, 427, _, _, 693, _, 146, 453, 321, 236, _, 444, 991, 1041, 
    841, 1234, 212, _, 536, _, _, 579, 1111, 565, 806, 2009, 937, 1934, 1172, 
    901, 481, 692, 239, 320, _, _, _, _, _, _, _, _, _, _, _, 2627, 1227, _, 
    2944, 5493, _, 458, 692, 145, _, _, _, _, _, _, _, _, _, _, 607, _, _, 
    1009, _, 858, 1174, _, 1086, _, 1142, _, 1326, 1371, 941, _, 1004, _, 
    295, _, 676, _, _, 275, 375, 857, 150, 163, 604, 621, 1412, _, 1729, _, 
    _, 570, 588, 361, 785, 924, _, 1773, _, 203, 316, 833, 142, 589, 208, 
    865, 1362, 7390, 306, 231, 2015, 2203, 2720, 786, 883, _, _, 2148, 187, 
    517, 2872, 583, 670, 1105, 447, _, 1304, 1191, _, 163, 311, 577, 274, 
    841, 1013, 784, 288, 668, _, 1609, 270, _, 944, 1199, 1398, _, 2240, 328, 
    _, _, _, _, 4484, _, 152, _, 983, _, 3882, 6523, 144, 355, 929, _, 2306, 
    704, 1423, 560, 720, 338, 1806, 505, 170, 439, 817, 2488, 761, 1452, 
    2689, _, _, _, _, _, 542, _, 985, 916, 1405, 916, _, _, _, _, _, _, _, 
    2843, 2518, 2485, 312, 2198, 1174, 2301, 796, _, 2365, 146, 240, 189, 
    178, 1710, 2531, 408, 2044, 221, _, _, 951, 844, 1204, _, _, _, _, _, 
    293, 1449, 780, 262, _, 705, 806, 165, 974, 460, 832, 1878, 490, 383, 
    377, 413, 415, _, _, 2525, 583, 186, 1712, 4339, 1542, 372, 338, 374, _, 
    _, _, _, _, _, 4550, 3967, 1187, 255, 792, 5022, 904, 745, 3115, 1471, 
    2835, 271, 1002, 874, _, 1146, _, 1202, _, 233, _, _, _, _, _, _, _, _, 
    1749, 2414, 4724, 4363, _, _, _, 6276, 6042, 3003, 11127, 9080, 12226, _, 
    _, _, _, 2271, 315, 388, _, 714, 1136, 577, _, _, 243, 1434, 7989, 8251, 
    _, 156, 172, 205, _, 469, 2007, _, _, 4301, 1356, 2338, 1856, 211, _, _, 
    _, _, 432, 1652, _, 614, 860, 782, 903, 966, _, 1427, 1308, 1287, 847, 
    1050, 1404, 1223, 562, 434, 579, 326, 247, 157, 139, _, 239, 267, _, _, 
    _, 2080, _, _, _, 2546, _, 2493, _, 206, _, _, _, _, 928, 964, _, 459, _, 
    2439, _, _, 3217, _, 1124, 520, _, 380, 1047, _, 1170, 1189, 1258, 898, 
    _, _, 1261, _, 1411, 2795, 3677, 2636, 328, 653, 816, 589, 876, 1833, 
    3210, 3935, _, 429, _, 573, 2050, 394, _, _, 2943, 1840, _, 1119, 1188, 
    _, _, _, 1639, 1738, 1815, 272, 990, _, _, _, _, _, _, 2967, 3820, 188, 
    592, 1163, 1628, 2645, 359, 398, 993, 844, 371, 464, 1683, 593, 4389, 
    727, _, 1780, 321, 295, 327, 212, 171, 1719, 486, _, _, _, 3818, 169, 
    1597, 141, 274, 771, 1147, _, _, 185, 205, 284, 344, 161, 603, 204, 333, 
    901, 134, 632, 1367, 435, _, _, 504, 336, _, 2147, 283, _, 269, 210, _, 
    628, 571, 854, 760, 235, 890, 1601, 1570, _, 2783, _, _, _, 2661, 2778, 
    2723, 5004, 4915, 747, _, 1002, 1046, 967, 1152, 383, 786, 222, _, 330, 
    720, 295, _, 1956, 507, 619, 164, _, 242, 539, 471, _, 151, 666, 3646, 
    3628, _, _, _, _, 1830, 2840, _, _, _, 2833, _, _, 2731, 4347, 1967, 505, 
    _, _, _, 783, _, _, 1049, _, 1135, 1319, _, 1507, _, _, 1133, _, _, 2636, 
    1782, _, 592, 1255, _, 3631, 1644, _, 1835, 1531, 1607, 1645, 2664, _, 
    22923, _, 660, 900, _, 692, 903, 1616, 724, 290, 362, 587, 482, 2226, 
    319, 364, _, 3010, 912, _, 674, 517, 1048, _, 1060, _, 1377, _, _, _, _, 
    _, _, _, 4513, 397, 1557, _, _, _, _, 184, 1073, 1806, 3151, 9010, _, 
    1401, _, 1993, 405, 367, 502, 353, 591, 561, 551, 1496, 969, 1122, 162, 
    383, 204, 1424, 523, 1917, _, _, _, _, _, _, _, 743, 685, 585, 244, 1468, 
    957, 248, _, 377, 261, _, _, 909, 835, 242, _, 459, 2802, 5232, 367, 
    1524, _, _, _, _, _, _, _, _, _, _, _, _, 9259, _, _, 1636, 1961, 2714, 
    3477, 1262, 1497, 1417, 1311, 1223, 313, 977, 759, 999, 1796, 928, 1334, 
    362, 250, 357, 434, 1176, 1905, 489, 265, 218, 4014, 437, 967, 266, 229, 
    332, 215, 382, 471, 1525, 448, 1052, 793, 490, 538, 256, 146, 258, 1521, 
    677, 287, 1193, 1986, _, _, _, _, _, _, _, _, _, _, 1295, 285, 445, 195, 
    354, 1746, 1254, _, 2429, 185, 853, 2220, 1292, 227, 153, 961, 711, 311, 
    153, 162, _, 140, _, _, _, _, _, _, _, _, _, _, _, _, _, 3732, 7208, _, 
    _, 4809, _, _, 3733, 2454, 2507, 993, 2642, 757, 159, 377, 1179, 179, 
    909, 245, 744, 536, 588, 369, 792, 916, 181, 782, 1164, 306, _, 815, 
    2058, _, _, _, _, _, _, 4036, _, 3104, _, 3261, 1348, 246, 629, _, 932, 
    1551, _, 2492, 2404, _, 974, _, 367, _, 601, _, 853, 13178, 2003, _, 
    8986, 7516, 8293, 8901, 1281, 1279, _, _, _, _, _, 1351, _, _, 1786, 
    1491, _, _, 1775, 1378, 704, 405, 562, 862, 283, 172, 526, 1132, 1028, 
    1134, 766, _, _, _, _, _, _, _, 1317, 1568, _, _, 406, 268, 228, 406, 
    309, 1086, _, 2256, 3003, 1049, 842, 792, _, 1030, _, 1135, _, _, 484, 
    812, _, 2265, 1871, _, _, _, _, 3466, 244, 478, 1450, 472, 606, 164, 269, 
    237, 172, 269, 170, 145, 220, 138, 183, 576, 403, 127, 124, 445, 1439, 
    1391, 264, 1264, _, _, _, 418, _, 279, _, 1155, 2176, 2277, 965, 1120, 
    2211, 1052, _, 2467, 193, 161, 302, 652, 576, _, 1904, 1563, 675, 542, 
    1113, 1393, 1259, 1417, _, _, _, _, _, _, _, _, _, _, 4744, 325, _, 267, 
    618, 2393, 413, _, 724, 1249, _, 3109, 3186, 356, 535, 880, 178, 350, 
    1127, _, 1779, 937, _, 402, 467, _, _, _, _, _, _, _, _, _, 3649, 350, 
    3658, 888, _, 445, _, 569, _, 638, 616, 842, _, 626, 842, 950, _, 174, 
    179, 505, 514, 747, 323, 645, 702, _, 1394, _, 263, 224, 725, 796, 5520, 
    _, 6332, _, _, _, _, _, 4249, _, 3220, _, _, _, _, _, _, _, _, _, 2459, 
    451, 168, 985, 1552, 184, _, 158, _, _, 794, 779, 757, 249, _, _, 678, 
    179, _, 451, 1871, _, _, 768, _, 1500, 1266, 975, 1228, 511, 967, 1227, 
    _, _, 3058, 2534, 1223, 4137, 2843, 557, 1651, 320, 869, _, 1788, _, _, 
    2024, 1718, 392, 246, 204, 519, 440, 320, 665, 387, 165, 2003, 434, 720, 
    1774, _, 4235, _, 2304, 1221, _, _, _, 1438, 1802, 1870, 683, 1106, 347, 
    568, 1139, 1574, 321, 1445, 1769, 1639, 1456, 741, 1374, 1237, 1269, 946, 
    _, 1630, 1640, 391, 941, 1737, _, _, _, _, _, _, _, _, 3697, 3549, _, 
    4347, _, _, _, 3683, 2906, 1341, 1362, _, 1375, 1331, 894, 195, 272, 618, 
    149, 853, 390, 511, 534, 972, 1054, _, _, 1253, 580, 2155, 193, _, 2411, 
    2392, _, _, 3279, 223, 1755, 2854, 2311, 2277, 2452, 429, 2704, 390, _, 
    417, 656, 187, 1193, 815, 385, 622, 166, 450, 650, 734, 650, 2141, 2299, 
    349, 373, 181, _, _, _, _, _, _, 3343, 2942, 2927, _, _, 532, 2868, _, _, 
    4209, 318, 347, 194, _, 528, _, _, 1634, _, 2781, 1175, _, 277, 724, _, 
    1264, _, 310, 1334, _, _, _, _, _, _, _, _, _, 2037, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, 3743, 2782, _, _, 859, _, 2953, _, 185, 266, 953, 
    2007, 3020, 1906, 1938, 1809, 3090, 226, 493, 2670, 4324, _, 5621, 689, 
    167, 773, 463, _, 758, _, _, 201, _, 206, 1010, 435, 507, 630, 733, 604, 
    412, 1282, 542, _, 706, 165, 218, 469, _, _, 933, 1176, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, 532, _, _, 756, 1683, 321, 571, 895, 1102, 
    1057, 1085, 1140, 1299, 1057, 251, 552, 305, 1221, 1541, 642, 994, _, 
    1394, _, _, _, _, 449, 4961, 350, 556, 251, 515, 127, 1059, _, 853, 1281, 
    198, 231, _, _, 159, 212, 750, _, 161, _, _, 928, 153, 486, 815, 195, 
    175, 739, _, 670, _, _, 795, 320, _, _, 1129, _, 6184, 365, 517, 401, 
    147, 236, 151, 198, 362, 700, 127, 352, 134, 336, 2860, 548, _, 657, 
    1923, 3848, _, 4693, 4102, 342, 201, 324, 441, 1786, 1351, 1186, 950, _, 
    _, 1246, _, 1330, 1419, _, 1484, 1275, 470, _, 914, _, 1063, 1276, 1601, 
    281, 643, 666, 983, 2324, 417, 268, 375, 283, 565, 936, 2543, 1997, 258, 
    479, 700, 880, 692, 558, 173, 154, 1042, 492, 1246, _, _, 646, 998, 1200, 
    590, 1773, 1084, _, _, _, 1474, 303, 224, 453, 407, 1112, 6573, 5218, 
    14145, 8984, 7879, 326, 181, 433, 382, 862, 129, _, 358, 329, 149, 229, 
    246, 1673, 1460, 411, 1391, 1185, 1186, _, 1077, _, _, _, 5121, 3181, 
    3366, 3517, _, 206, _, 1185, _, 524, 405, 455, _, 966, 575, 3912, 1182, 
    3082, 5030, 1962, 638, 321, _, _, _, 2555, _, _, 2595, _, _, _, _, 3439, 
    532, 1000, 1127, _, 213, 906, 156, 220, 479, _, _, 1086, 5804, 1085, 
    1147, 3809, 289, 11441, 7691, _, 9657, 1535, 302, 174, 219, 2473, 5868, 
    5764, 206, 178, 340, 895, 1071, 1325, 1417, 1276, 937, 1429, 1525, 1388, 
    _, _, _, _, 1479, 216, 883, 501, 184, 147, _, _, _, _, 2722, 2220, 2239, 
    869, 465, 1173, 2647, 799, 161, 199, 255, _, 3872, 590, 399, 446, 633, 
    556, 150, 528, 505, _, 451, 443, 520, _, 806, _, 890, 932, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, 3562, _, _, _, 276, _, 708, _, 764, 584, _, 1699, 
    475, 2298, 144, 1097, 626, 524, 233, 1008, 247, 618, 161, 274, 151, 916, 
    142, 838, 225, 599, 777, _, _, _, _, 13262, _, 415, _, 1884, 2719, 428, 
    329, 442, 139, 152, 1813, 2115, 140, 158, 182, 163, 2900, 5105, 152, 159, 
    742, 534, 186, 934, _, _, _, _, _, _, _, _, 391, _, 1009, _, 1074, 1319, 
    _, _, 1507, 1515, 494, _, _, 618, 716, _, 644, _, 2088, 326, 510, _, 576, 
    _, 201, 241, 695, 1388, 1787, _, 2752, _, 3475, _, _, 707, 999, 1086, _, 
    _, 1429, _, _, 1214, 3189, _, 592, _, _, 767, 140, _, _, 944, 208, 411, 
    _, 2609, _, _, 1947, 6561, 9141, 1046, 1277, _, _, _, 1215, 2756, _, 
    1640, 2800, _, 332, 213, 297, 198, _, 259, _, _, _, 578, 567, _, 820, 
    512, 1743, 7125, _, 7240, 1130, _, _, _, 1781, 1574, _, _, 1777, _, _, 
    172, _, 554, _, 428, _, 2196, 486, 725, 1386, 1116, 451, 875, 1704, 1764, 
    1500, 1180, 984, _, _, _, _, 5354, 4770, _, 1748, 2187, 807, _, 1916, _, 
    186, _, 210, 2553, 3051, 3714, 6722, 3739, 237, 928, 1200, 160, _, 742, 
    1225, _, _, _, 1556, _, _, 1572, 463, 677, 536, 487, _, _, _, _, _, _, 
    436, _, 1058, 1128, 1350, _, _, 1118, 1207, 1355, 938, 1299, 1434, 1174, 
    725, 985, _, 761, _, 1221, _, _, 1713, _, _, 1873, 2020, 2361, 1307, _, 
    1457, 1411, 138, 354, 484, 677, _, 1072, 158, _, _, _, _, _, 2080, _, 
    1592, _, 290, 187, 170, 2346, 2884, 753, 724, 906, 1023, 581, _, 2663, 
    2478, _, 1026, 3834, 5742, 7305, 6323, 1232, 7156, 448, 469, 2237, 400, 
    542, 467, 643, 2172, 324, 724, 1010, 671, 571, 247, 365, 1153, _, 1726, 
    1351, 230, 245, 973, 2151, 1297, _, _, _, _, 2506, _, _, 4606, 3934, 
    3985, 568, 1146, 551, 1106, 504, _, _, _, _, 1600, 1583, _, 673, 626, 
    462, 141, 867, 528, 397, 148, 293, 768, 528, 115, 115, 163, 281, 246, 
    190, 446, 822, 223, 350, 832, 582, 350, 363, 402, 260, 4278, 3825, _, 
    278, 535, 1110, 1699, 269, _, 1884, 246, 645, 567, 665, 1030, 926, 917, 
    1439, 1181, 2952, 232, 679, 1113, 947, _, 1577, 954, _, 1124, 265, _, _, 
    5186, 941, 1689, 798, 700, 467, 1123, 276, _, 334, 461, 416, 985, 1469, 
    1043, 152, 308, 607, _, 3083, _, _, _, 7668, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, 13632, 28013, _, 3273, 3997, 1079, 423, 497, 856, 220, 
    956, 213, 318, _, 212, 382, _, _, 185, _, 367, _, 439, 1520, _, 2860, 
    2023, 919, 407, _, _, 900, _, 2165, _, _, _, _, 3535, 1507, 1464, 883, 
    1391, 1609, 2419, _, 1016, _, 271, _, 495, 557, 190, 363, 399, _, 434, 
    332, 934, 4928, 3704, 661, _, _, 2156, 698, 1805, 236, 150, 3046, 3677, 
    512, 266, 833, 505, 748, 761, 143, 402, 376, 655, 763, 151, 125, 387, 
    480, 186, 203, 502, 1070, 177, 212, 510, 1504, 8706, 347, 1332, 3357, 
    581, 768, _, 447, 567, 3798, 1839, _, 880, 731, _, _, _, _, 1163, _, _, 
    1407, _, _, 1399, _, _, 1477, _, 254, _, _, _, _, _, 439, 1240, _, 352, 
    _, _, _, 145, 138, 305, 3595, 1123, _, 1595, 392, 828, 916, 1067, 826, _, 
    _, 3219, _, _, _, _, 3790, 3290, _, 2228, 2107, _, 456, 501, _, 1150, 
    1091, 885, 275, 478, 708, 1070, 1176, 1249, 1189, _, _, 1535, 2119, _, _, 
    2653, 2656, 9380, 8330, 6934, 302, 737, 523, 457, 926, _, _, _, 1065, 
    305, 261, 2082, 395, 814, 788, 712, 935, 178, 519, 521, 155, 1020, 455, 
    1827, 406, 641, 781, 748, 1003, 706, 700, 715, 546, _, _, 1342, 1314, _, 
    _, 1451, 996, 1093, 1882, 162, _, 1864, 1647, _, 927, _, _, _, 222, 269, 
    677, 1923, 2188, 575, 241, 375, 733, 1323, 620, 773, 412, 273, 382, 2521, 
    1254, 304, 581, _, 1396, _, 2153, 1938, _, _, _, 1680, _, 593, _, _, 357, 
    730, 385, _, 464, _, 397, _, _, _, _, _, _, _, 1615, _, 266, _, 584, 586, 
    271, 525, 786, 499, 2403, 2090, 101738, 163345, 167422, 1162, 971, 497, 
    821, 734, _, 1085, 1314, 1778, 2721, _, 2478, 1880, _, 553, 1082, 1197, 
    1537, _, _, _, _, _, _, _, _, _, _, 256, 579, 801, 758, 934, 1106, 379, 
    216, 141, 238, 150, 217, 307, 168, 997, 157, 169, 399, 241, 260, 239, 
    418, 190, 815, 860, _, _, 618, 352, 359, _, 537, 794, 701, _, 1150, _, _, 
    _, 1815, 1974, _, _, 2097, 1046, _, 216, 138, _, 618, 1006, 1276, 204, 
    390, 1661, 928, 217, 736, 164, 318, 535, 842, 160, 551, 668, 272, 230, _, 
    204, 519, 210, 796, 538, 190, 384, _, 221, 298, 876, 853, 412, 495, 488, 
    3680, _, 4752, 5472, 993, _, _, 1724, _, _, _, _, _, _, _, _, 2095, 338, 
    389, 644, _, _, 636, 587, 468, 1164, 847, 263, 399, 173, 432, 1629, 794, 
    _, 986, 776, 495, _, _, 358, _, _, 630, 386, 588, 1194, 431, 794, 1015, 
    _, _, _, _, _, _, _, _, 4019, _, _, _, 972, 1582, 796, 687, 625, 1149, 
    269, 237, 220, 204, 245, 501, 405, 382, 346, 252, 868, 518, 180, 676, _, 
    644, 284, 275, 1482, _, 1858, _, 1452, 158, 219, 1700, 1621, 2062, 3263, 
    1126, 1235, _, 173, _, 816, 284, 2197, 1446, 558, 561, 6256, 351, 4361, 
    4381, 620, 667, 2118, 735, 480, 1136, 2422, 254, 417, 122, 346, 186, 
    1096, 869, 602, 169, 778, 780, 887, _, 1230, 906, 474, _, _, _, _, _, _, 
    _, 3487, 3487, 655, _, 2315, 2651, 3879, 1318, 2168, 2191, 2201, 987, 
    325, 858, 535, 160, 1330, 11142, 386, 1055, 613, 807, 980, 2444, 2076, 
    1011, 1591, 2102, 3150, 2855, 166, 192, 2448, 2871, _, _, 2734, 2475, 
    1797, 254, 349, 783, 952, 262, 284, 279, 286, 361, 735, 948, 9518, 2846, 
    1791, 4450, _, 4643, 921, 306, 268, 891, _, _, _, _, 11659, _, _, _, 
    1033, 657, 562, _, 569, 239, 216, 381, 489, 273, 527, _, 2127, 2162, 290, 
    _, 298, 577, 1138, 1521, 3411, 4857, 3018, 4388, 214, 1685, 542, 354, 
    413, 215, 214, _, _, 567, 255, 632, 804, 822, _, 878, 921, 215, 808, 
    1317, _, _, _, _, _, 2304, _, _, 222, 298, 363, 315, 301, _, _, _, 1973, 
    516, 634, _, _, 1180, 2959, 3208, 5455, 2850, 876, 2065, 2770, 627, 825, 
    1135, 1218, 1297, 1490, 1044, _, 711, _, 3161, _, 2272, 578, 1031, 856, 
    825, _, _, 442, _, _, _, _, _, _, 421, 645, 421, 196, 493, 362, 441, 
    1320, 203, 321, 280, _, _, 938, 189, 1461, 1304, 826, 1019, 4516, _, 
    5363, 2277, 1106, 1377, _, _, _, _, 772, 2550, _, 2906, 1147, _, 507, _, 
    _, _, _, 8543, 10768, _, _, 7795, _, 2139, _, _, 2243, 316, 443, _, 484, 
    _, 747, 337, _, 1060, 1064, 1142, 1304, 1431, 1091, 681, 286, 791, 973, 
    _, 845, 667, 1042, _, 377, 159, 122, 857, 182, 1943, 151, 256, 325, _, 
    201, 191, 537, 537, 1261, 2221, _, 619, 974, 1053, 4662, 2003, _, _, 
    6319, _, _, 905, 146, 520, 770, _, _, _, _, 266, _, _, 1753, 1512, 875, 
    944, 591, 616, 1173, 331, _, 386, 392, 469, 437, 1768, 406, 5634, _, 
    7697, _, 369, 1022, 1223, 1400, 2938, _, 2827, 3761, 645, _, 2376, 1200, 
    1144, 1372, 1236, _, _, 1901, 1208, 616, 808, 1489, 483, 1185, 1333, 
    1320, 710, 1941, _, 726, 783, 828, 278, 934, 873, 370, 2434, _, 2176, _, 
    _, _, 249, 186, 154, 172, 185, 1827, 3367, 2554, 1496, 730, _, 2123, 207, 
    _, 213, _, _, _, 210, _, 388, _, 283, 1217, 2981, 1045, 1374, _, _, _, _, 
    _, _, _, 7084, 685, _, _, 3232, 2721, 650, 153, 193, 913, 741, 691, 1484, 
    3601, 2754, 1042, 1424, 885, 393, 215, 173, 1236, 1260, 1596, 1939, 244, 
    _, _, _, _, 2714, 2147, 1281, 1790, 894, 707, _, 998, _, 1757, 3145, _, 
    730, 857, 961, 858, 246, _, 1164, _, _, _, _, _, _, _, 1397, _, _, 313, 
    1188, _, 2347, 580, 238, 309, 3048, 758, 759, 551, 318, 255, 260, 1907, 
    1415, 448, 863, 871, _, _, _, _, _, _, 1184, _, 329, 478, 1874, 879, 234, 
    362, _, 144, 724, 874, 495, _, 2772, 1804, 2002, _, 1948, 1746, 1525, 
    355, 769, 317, 396, 1687, 197, 363, 375, 414, 687, 949, 2570, 2590, 2921, 
    500, 1270, _, 748, 342, _, _, _, 1513, _, 1371, 256, 212, 179, 1916, 578, 
    1340, 288, _, 445, 1161, 909, _, 1601, _, 1733, _, 384, _, _, 205, _, 
    482, _, 379, 3488, _, 260, 258, 831, 1278, 1262, 439, 306, 719, 1000, 
    313, 229, 1562, 2169, 1443, 2031, 3586, 1164, 221, 231, 974, 1137, 2035, 
    267, 529, 202, 1131, 1387, 227, 1182, 174, 815, 853, 1051, 1140, 190, 
    538, 154, 671, 190, 462, 519, 239, 2084, 1748, 633, 621, 532, 417 ;

 instrument_location = _ ;

 instrument_pressure = _ ;

 instrument_tag = _ ;

 lat = 59.0913, 59.0941, 59.0955, 59.0995, 59.1, 59.0973, 59.1098, 59.1222, 
    59.1901, 59.1804, 59.1779, 59.183, 59.1832, 59.1929, 59.2031, 59.1965, 
    59.1924, 59.1859, 59.1959, 59.1918, 59.1893, 59.1925, 59.1861, 59.1899, 
    59.1933, 59.1869, 59.1814, 59.179, 59.185, 59.1874, 59.1885, 59.1896, 
    59.1896, 59.1809, 59.1846, 59.1822, 59.1844, 59.1776, 59.1571, 59.1543, 
    59.1355, 59.1072, 59.0952, 59.095, 59.0931, 59.0923, 59.0936, 59.0937, 
    59.0904, 59.0938, 59.0959, 59.0954, 59.1037, 59.113, 59.1225, 59.1351, 
    59.1466, 59.1561, 59.1627, 59.1721, 59.0942, 59.179, 59.1892, 59.1046, 
    59.1885, 59.1571, 59.1859, 59.185, 59.1927, 59.1979, 59.2009, 59.2143, 
    59.2056, 59.2147, 59.2226, 59.1864, 59.2044, 59.1968, 59.2012, 59.2169, 
    59.2134, 59.222, 59.2139, 59.2203, 59.1907, 59.1987, 59.2236, 59.2065, 
    59.2193, 59.2251, 59.2235, 59.2345, 59.2225, 59.2159, 59.2107, 59.211, 
    59.211, 59.1943, 59.1935, 59.1926, 59.1869, 59.1873, 59.1892, 59.1809, 
    59.1923, 59.1799, 59.1822, 59.1877, 59.1846, 59.1847, 59.1882, 59.1969, 
    59.1969, 59.1927, 59.2141, 59.194, 59.1874, 59.1926, 59.1925, 59.1931, 
    59.1984, 59.1845, 59.1986, 59.1978, 59.198, 59.1951, 59.1927, 59.1736, 
    59.1789, 59.1781, 59.1784, 59.1839, 59.1817, 59.1817, 59.1774, 59.1783, 
    59.1783, 59.1714, 59.1687, 59.1705, 59.1682, 59.181, 59.1799, 59.1803, 
    59.18, 59.1854, 59.169, 59.1839, 59.1982, 59.1994, 59.1921, 59.2002, 
    59.2003, 59.2019, 59.1979, 59.1978, 59.1978, 59.1977, 59.1975, 59.1943, 
    59.1931, 59.1938, 59.193, 59.1936, 59.1934, 59.1939, 59.1941, 59.1908, 
    59.1966, 59.1982, 59.1937, 59.1968, 59.1939, 59.199, 59.1964, 59.1884, 
    59.176, 59.1935, 59.1766, 59.1768, 59.1821, 59.1935, 59.1934, 59.1965, 
    59.1922, 59.1972, 59.1888, 59.1907, 59.1955, 59.195, 59.1947, 59.1963, 
    59.1956, 59.1937, 59.1937, 59.1894, 59.1853, 59.1785, 59.1889, 59.1571, 
    59.1166, 59.1042, 59.0999, 59.1201, 59.1177, 59.1216, 59.1294, 59.1183, 
    59.1614, 59.1552, 59.1546, 59.1583, 59.1577, 59.1568, 59.1743, 59.1527, 
    59.1618, 59.1725, 59.1711, 59.175, 59.1745, 59.174, 59.172, 59.1729, 
    59.1761, 59.1762, 59.1695, 59.1884, 59.1953, 59.1954, 59.2051, 59.1835, 
    59.2058, 59.2061, 59.1986, 59.2027, 59.209, 59.2062, 59.2113, 59.2097, 
    59.2089, 59.2087, 59.2104, 59.2178, 59.2103, 59.2113, 59.2097, 59.2153, 
    59.2075, 59.2077, 59.2147, 59.2136, 59.2108, 59.2077, 59.2073, 59.1543, 
    59.1243, 59.113, 59.1192, 59.1183, 59.1145, 59.1183, 59.1147, 59.1222, 
    59.1264, 59.2104, 59.1484, 59.1477, 59.1657, 59.1688, 59.1634, 59.1634, 
    59.1607, 59.1586, 59.1619, 59.1511, 59.1168, 59.0951, 59.1004, 59.0945, 
    59.0863, 59.0951, 59.1144, 59.0951, 59.0948, 59.0934, 59.0932, 59.0961, 
    59.0937, 59.0958, 59.0946, 59.0933, 59.0981, 59.0943, 59.0984, 59.1038, 
    59.1184, 59.1042, 59.1612, 59.1315, 59.1249, 59.1164, 59.1214, 59.1152, 
    59.109, 59.1107, 59.1163, 59.1237, 59.1162, 59.1097, 59.1101, 59.1203, 
    59.105, 59.1113, 59.1128, 59.1144, 59.1182, 59.1264, 59.1354, 59.0093, 
    59.12, 59.1137, 59.1168, 59.1153, 59.1145, 59.1264, 59.1234, 59.1261, 
    59.1191, 59.1251, 59.1267, 59.1262, 59.1215, 59.1217, 59.1213, 59.1249, 
    59.1155, 59.1191, 59.1214, 59.1293, 59.0916, 59.1234, 59.1165, 59.0935, 
    59.0945, 59.1154, 59.1084, 59.1099, 59.1163, 59.1223, 59.1297, 59.1295, 
    59.0951, 59.0994, 59.0971, 59.0927, 59.0916, 59.0946, 59.0935, 59.0935, 
    59.0926, 59.1001, 59.0999, 59.094, 59.0926, 59.0939, 59.0939, 59.0968, 
    59.0938, 59.0953, 59.0986, 59.0962, 59.0949, 59.0972, 59.0961, 59.0954, 
    59.0833, 59.0926, 59.0993, 59.0949, 59.097, 59.0899, 59.0871, 59.0984, 
    59.1393, 59.1457, 59.1467, 59.1673, 59.1673, 59.1561, 59.146, 59.1482, 
    59.1409, 59.1385, 59.137, 59.1275, 59.1222, 59.1109, 59.1098, 59.0902, 
    59.1013, 59.1106, 59.0999, 59.1055, 59.1061, 59.1058, 59.109, 59.1069, 
    59.1063, 59.1071, 59.1088, 59.107, 59.1069, 59.1045, 59.1073, 59.1166, 
    59.086, 59.098, 59.1071, 59.1101, 59.1542, 59.1614, 59.1545, 59.1519, 
    59.178, 59.1868, 59.1833, 59.1885, 59.1941, 59.1971, 59.0324, 59.1997, 
    59.2218, 59.2278, 59.2103, 59.1925, 59.201, 59.1983, 59.1959, 59.1882, 
    59.182, 59.1936, 59.1753, 59.175, 59.1759, 59.1624, 59.1587, 59.1593, 
    59.1453, 59.1269, 59.1253, 59.1159, 59.1258, 59.1248, 59.1165, 59.1144, 
    59.1226, 59.1193, 59.0913, 59.116, 59.1164, 59.1305, 59.096, 59.1119, 
    59.1132, 59.1038, 59.1591, 59.1598, 59.1642, 59.1629, 59.1623, 59.1613, 
    59.1612, 59.2172, 59.1576, 59.1836, 59.1585, 59.1704, 59.1431, 59.157, 
    59.1555, 59.1755, 59.1756, 59.1761, 59.1752, 59.1478, 59.1328, 59.1158, 
    59.1199, 59.1204, 59.1281, 58.9966, 59.1301, 59.1294, 59.1281, 59.127, 
    59.0762, 59.0944, 59.0876, 59.0905, 59.081, 59.0926, 59.0962, 59.1085, 
    59.0661, 59.0692, 59.0969, 59.1117, 59.1025, 59.0721, 59.1012, 59.1132, 
    59.1148, 59.117, 59.1206, 59.1201, 59.1297, 59.1178, 59.1167, 59.1239, 
    59.1169, 59.1155, 59.114, 59.1152, 59.1159, 59.1171, 59.1194, 59.119, 
    59.1189, 59.1186, 59.1189, 59.1187, 59.1192, 59.1186, 59.1211, 59.1145, 
    59.1196, 59.122, 59.1196, 59.0987, 59.0951, 59.0974, 59.099, 59.0902, 
    59.0919, 59.0999, 59.0992, 59.1013, 59.0997, 59.1042, 59.1002, 59.1074, 
    59.0974, 59.0986, 59.1043, 59.1009, 59.1069, 59.0961, 59.0959, 59.1002, 
    59.0959, 59.0967, 59.0979, 59.0954, 59.0919, 59.0928, 59.0967, 59.101, 
    59.096, 59.1121, 59.1181, 59.1187, 59.1247, 59.1246, 59.125, 59.1141, 
    59.1098, 59.1238, 59.1359, 59.1363, 59.1358, 59.1438, 59.2077, 59.2076, 
    59.2021, 59.1947, 59.1919, 59.1838, 59.0459, 59.1223, 59.1459, 59.1518, 
    59.1446, 59.1526, 59.1136, 59.1196, 59.1242, 59.1287, 59.1026, 59.0994, 
    59.0978, 59.1055, 59.1111, 59.1133, 59.1045, 59.1019, 59.0987, 59.1071, 
    59.0892, 59.0858, 59.0874, 59.0959, 59.0988, 59.0952, 59.0794, 59.0845, 
    59.1257, 59.1574, 59.1492, 59.1645, 59.1849, 59.2021, 59.1965, 59.1964, 
    59.197, 59.2055, 59.2375, 59.1928, 59.1937, 59.196, 59.2176, 59.207, 
    59.2068, 59.2093, 59.1745, 59.1835, 59.1856, 59.1753, 59.1731, 59.2181, 
    59.22, 59.2212, 59.2217, 59.2243, 59.207, 59.2294, 59.2213, 59.219, 
    59.2172, 59.2199, 59.2239, 59.2217, 59.2179, 59.2258, 59.2175, 59.2193, 
    59.2224, 59.2247, 59.2184, 59.2146, 59.2138, 59.2122, 59.2157, 59.1799, 
    59.1855, 59.1883, 59.183, 59.1827, 59.1826, 59.1847, 59.1944, 59.1881, 
    59.2029, 59.2016, 59.2009, 59.1985, 59.1985, 59.196, 59.1976, 59.1993, 
    59.1928, 59.1625, 59.1876, 59.1674, 59.1753, 59.1889, 59.1998, 59.2046, 
    59.1793, 59.1941, 59.1941, 59.2006, 59.196, 59.1997, 59.2007, 59.1664, 
    59.1998, 59.1509, 59.1775, 59.1519, 59.1768, 59.1517, 59.1572, 59.1677, 
    59.1739, 59.1736, 59.1748, 59.1625, 59.1855, 59.1821, 59.182, 59.1878, 
    59.1886, 59.1951, 59.2083, 59.2189, 59.2198, 59.2271, 59.2216, 59.226, 
    59.2187, 59.2186, 59.2185, 59.2188, 59.2438, 59.2363, 59.218, 59.2263, 
    59.2206, 59.2178, 59.2198, 59.219, 59.2206, 59.2184, 59.2201, 59.2167, 
    59.2153, 59.2493, 59.2192, 59.2194, 59.2177, 59.2195, 59.2178, 59.2169, 
    59.2184, 59.2204, 59.2268, 59.216, 59.2186, 59.2187, 59.2226, 59.2188, 
    59.1898, 59.1828, 59.1835, 59.1908, 59.1923, 59.182, 59.345, 59.2235, 
    59.1494, 59.1426, 59.1323, 59.1441, 59.1076, 59.0902, 59.0993, 59.0982, 
    59.1434, 59.0949, 59.094, 59.0981, 59.0971, 59.0962, 59.095, 59.0866, 
    59.0936, 59.0843, 59.0927, 59.0942, 59.0943, 59.0801, 59.0926, 59.1334, 
    59.1392, 59.1427, 59.1615, 59.1889, 59.1847, 59.1825, 59.2479, 59.2454, 
    59.0627, 59.073, 59.2178, 59.2154, 59.2066, 59.2186, 59.2139, 59.1994, 
    59.2036, 59.1943, 59.1926, 59.1725, 59.1719, 59.1792, 59.1952, 59.1928, 
    59.2031, 59.2082, 59.2083, 59.2085, 59.1767, 59.1763, 59.2073, 59.176, 
    59.2059, 59.1439, 59.1797, 59.1943, 59.1926, 59.1893, 59.1873, 59.1916, 
    59.1918, 59.1928, 59.193, 59.1937, 59.1957, 59.1847, 59.197, 59.1983, 
    59.2435, 59.2609, 59.2738, 59.2738, 59.2826, 59.27, 59.2698, 59.2961, 
    59.3033, 59.2579, 59.2593, 59.2315, 59.2004, 59.2072, 59.1976, 59.1971, 
    59.1975, 59.2774, 59.192, 59.1892, 59.173, 59.1912, 59.1958, 59.1925, 
    59.187, 59.2043, 59.2039, 59.2041, 59.1982, 59.202, 59.202, 59.2038, 
    59.2032, 59.2027, 59.2046, 59.2022, 59.1653, 59.1629, 59.1838, 59.1776, 
    59.1783, 59.172, 59.1548, 59.1731, 59.1785, 59.1814, 59.1636, 59.1637, 
    59.1784, 59.1896, 59.1796, 59.1758, 59.1914, 59.1821, 59.1833, 59.1886, 
    59.1228, 59.102, 59.1269, 59.1349, 59.1821, 59.1809, 59.1828, 59.191, 
    59.1839, 59.1749, 59.2298, 59.1941, 59.1884, 59.1885, 59.1842, 59.1812, 
    59.1924, 59.191, 59.1956, 59.1937, 59.1916, 59.1967, 59.1977, 59.1988, 
    59.1747, 59.1844, 59.186, 59.1606, 59.1589, 59.1567, 59.1545, 59.1744, 
    59.1825, 59.1543, 59.1712, 59.1694, 59.1651, 59.1655, 59.1793, 59.177, 
    59.1831, 59.1135, 59.1891, 59.1898, 59.1935, 59.1955, 59.1936, 59.1908, 
    59.1973, 59.1969, 59.1934, 59.1799, 59.1906, 59.1861, 59.1894, 59.1904, 
    59.1928, 59.1864, 59.1895, 59.1896, 59.1893, 59.1886, 59.1792, 59.1926, 
    59.1818, 59.1669, 59.1872, 59.1031, 59.125, 59.1168, 59.1168, 59.1162, 
    59.1159, 59.1162, 59.1252, 59.1251, 59.1295, 59.1277, 59.1182, 59.1059, 
    59.0949, 59.0874, 59.0872, 59.0873, 59.0978, 59.0974, 59.0971, 59.0951, 
    59.0957, 59.093, 59.095, 59.0952, 59.0962, 59.0961, 59.0961, 59.0938, 
    59.0942, 59.097, 59.1002, 59.0925, 59.1094, 59.0966, 59.0952, 59.0886, 
    59.0886, 59.0918, 59.1175, 59.1176, 59.1295, 59.1147, 59.1101, 59.0931, 
    59.1115, 59.1189, 59.1189, 59.1309, 59.142, 59.129, 59.1292, 59.1215, 
    59.1152, 59.1121, 59.1198, 59.1112, 59.1102, 59.1107, 59.1327, 59.1328, 
    59.1638, 59.1641, 59.1847, 59.1921, 59.1931, 59.1929, 59.2, 59.1926, 
    59.202, 59.2079, 59.206, 59.201, 59.195, 59.2006, 59.136, 59.1417, 
    59.1409, 59.1762, 59.1457, 59.186, 59.1912, 59.1916, 59.2079, 59.1893, 
    59.1805, 59.1853, 59.1812, 59.1838, 59.2026, 59.1951, 59.2072, 59.195, 
    59.1901, 59.1975, 59.2019, 59.1847, 59.2177, 59.2179, 59.2233, 59.1987, 
    59.1629, 59.1979, 59.1979, 59.1926, 59.1959, 59.1964, 59.179, 59.1793, 
    59.1905, 59.1912, 59.1914, 59.1912, 59.201, 59.1959, 59.1927, 59.1952, 
    59.1971, 59.1951, 59.1912, 59.1924, 59.186, 59.1922, 59.1946, 59.1922, 
    59.1934, 59.1922, 59.1895, 59.192, 59.1969, 59.1915, 59.1797, 59.1779, 
    59.1712, 59.1631, 59.1564, 59.2702, 59.1594, 59.1656, 59.1717, 59.1793, 
    59.1742, 59.1729, 59.167, 59.1685, 59.1758, 59.1795, 59.1824, 59.1822, 
    59.1824, 59.18, 59.1768, 59.184, 59.1826, 59.1757, 59.1756, 59.1669, 
    59.1711, 59.1703, 59.1749, 59.1841, 59.19, 59.1732, 59.1909, 59.1744, 
    59.1976, 59.1969, 59.1907, 59.19, 59.19, 59.1946, 59.194, 59.1946, 
    59.1997, 59.1948, 59.1975, 59.1953, 59.1978, 59.1931, 59.1951, 59.1968, 
    59.1929, 59.1996, 59.195, 59.1954, 59.1969, 59.1946, 59.1969, 59.1954, 
    59.1953, 59.1938, 59.1946, 59.1996, 59.1945, 59.1945, 59.1908, 59.1863, 
    59.1873, 59.1942, 59.1851, 59.1951, 59.1956, 59.1806, 59.2131, 59.2054, 
    59.1799, 59.1824, 59.1822, 59.1821, 59.1757, 59.1722, 59.1752, 59.1881, 
    59.2278, 59.2372, 59.156, 59.1569, 59.1628, 59.1843, 59.1928, 59.1912, 
    59.1922, 59.1945, 59.1946, 59.1933, 59.1959, 59.1917, 59.1956, 59.1967, 
    59.1929, 59.193, 59.1975, 59.1923, 59.1828, 59.181, 59.174, 59.1864, 
    59.1834, 59.1825, 59.1938, 59.2041, 59.149, 59.1332, 59.2327, 59.1535, 
    59.139, 59.1841, 59.1806, 59.1446, 59.1181, 59.1065, 59.194, 59.1464, 
    59.1858, 59.1951, 59.2059, 59.2111, 59.1933, 59.2445, 59.1905, 59.2015, 
    59.1838, 59.1686, 59.1626, 59.1313, 59.1791, 59.1202, 59.1184, 59.1072, 
    59.0969, 59.0975, 59.1224, 59.0775, 59.1151, 59.1301, 59.0979, 59.0919, 
    59.0944, 59.094, 59.0924, 59.092, 59.0917, 59.0921, 59.0886, 59.0966, 
    59.1005, 59.0841, 59.1158, 59.123, 59.1193, 59.125, 59.1292, 59.181, 
    59.1811, 59.181, 59.181, 59.181, 59.1542, 59.1881, 59.1963, 59.1922, 
    59.1923, 59.1912, 59.1907, 59.1898, 59.1914, 59.1996, 59.2111, 59.2036, 
    59.1819, 59.1805, 59.182, 59.1783, 59.1782, 59.1701, 59.1704, 59.1708, 
    59.1703, 59.1774, 59.1771, 59.1748, 59.1761, 59.1759, 59.1742, 59.1752, 
    59.1734, 59.1754, 59.1737, 59.1767, 59.1608, 59.1745, 59.1792, 59.1764, 
    59.1836, 59.197, 59.2084, 59.1968, 59.196, 59.1973, 59.1708, 59.1385, 
    59.1076, 59.0894, 59.0906, 59.095, 59.0961, 59.0901, 59.0974, 59.0964, 
    59.0963, 59.0978, 59.0985, 59.094, 59.0965, 59.0962, 59.0947, 59.0972, 
    59.0939, 59.0947, 59.0971, 59.0853, 59.085, 59.0749, 59.1535, 59.1915, 
    59.1892, 59.1753, 59.1709, 59.1937, 59.171, 59.1751, 59.1891, 59.1939, 
    59.2023, 59.1962, 59.1905, 59.1926, 59.1942, 59.1925, 59.1926, 59.1911, 
    59.1991, 59.2103, 59.2099, 59.2067, 59.2018, 59.2016, 59.2246, 59.2052, 
    59.1968, 59.1984, 59.1945, 59.1905, 59.1984, 59.2005, 59.2043, 59.1961, 
    59.2101, 59.2177, 59.2256, 59.2305, 59.228, 59.2244, 59.2174, 59.2182, 
    59.2179, 59.2161, 59.199, 59.1958, 59.194, 59.1935, 59.1736, 59.1723, 
    59.1922, 59.1794, 59.1766, 59.1844, 59.191, 59.1873, 59.1892, 59.1861, 
    59.1902, 59.1831, 59.1783, 59.1808, 59.1843, 59.1862, 59.1881, 59.1926, 
    59.1784, 59.1738, 59.1614, 59.1589, 59.1582, 59.1532, 59.1381, 59.137, 
    59.1294, 59.1206, 59.093, 59.0926, 59.1078, 59.0977, 59.0914, 59.0896, 
    59.0801, 59.0914, 59.1025, 59.096, 59.0973, 59.1002, 59.0982, 59.1098, 
    59.1082, 59.0999, 59.0822, 59.0766, 59.0951, 59.0899, 59.0867, 59.0979, 
    59.0979, 59.095, 59.0951, 59.0979, 59.0972, 59.0922, 59.0924, 59.1271, 
    59.1337, 59.2174, 59.1966, 59.2268, 59.2359, 59.2381, 59.2374, 59.2419, 
    59.235, 59.1792, 59.1717, 59.1865, 59.2234, 59.2258, 59.2186, 59.1964, 
    59.21, 59.2225, 59.2149, 59.2001, 59.2002, 59.2173, 59.2234, 59.2218, 
    59.2097, 59.2173, 59.2221, 59.2204, 59.2273, 59.2105, 59.2086, 59.2031, 
    59.204, 59.2019, 59.2056, 59.2036, 59.1976, 59.1921, 59.1894, 59.1935, 
    59.1932, 59.1879, 59.1673, 59.2186, 59.2091, 59.1977, 59.1623, 59.1624, 
    59.155, 59.1456, 59.1573, 59.1437, 59.1476, 59.149, 59.2194, 59.2188, 
    59.2188, 59.2259, 59.2238, 59.2131, 59.1768, 59.16, 59.1557, 59.151, 
    59.1461, 59.1502, 59.1485, 59.1342, 59.1283, 59.1307, 59.0932, 59.0907, 
    59.0927, 59.093, 59.0961, 59.0939, 59.0946, 59.1176, 59.1191, 59.113, 
    59.106, 59.0984, 59.1131, 59.1282, 59.1214, 59.105, 59.0943, 59.0961, 
    59.0778, 59.119, 59.1643, 59.1832, 59.1748, 59.157, 59.1503, 59.1446, 
    59.1502, 59.1212, 59.1147, 59.1087, 59.1128, 59.1211, 59.1315, 59.1323, 
    59.1119, 59.0999, 59.0961, 59.0936, 59.0906, 59.085, 59.0979, 59.0891, 
    59.1057, 59.112, 59.1166, 59.108, 59.136, 59.2041, 59.1853, 59.1848, 
    59.1042, 59.0956, 59.0949, 59.095, 59.095, 59.0954, 59.0949, 59.0994, 
    59.095, 59.1014, 59.0949, 59.0998, 59.0954, 59.0934, 59.0965, 59.1006, 
    59.0961, 59.106, 59.096, 59.0946, 59.094, 59.094, 59.094, 59.0962, 
    59.0934, 59.0952, 59.0933, 59.0958, 59.0964, 59.1622, 59.1633, 59.0902, 
    59.0914, 59.1078, 59.1092, 59.7264, 59.2752, 59.205, 59.2288, 59.215, 
    59.2238, 59.2063, 59.2101, 59.2152, 59.2103, 59.2076, 59.2106, 59.21, 
    59.2277, 59.2115, 59.2118, 59.2116, 59.2057, 59.2096, 59.2094, 59.2033, 
    59.2092, 59.2091, 59.2084, 59.2154, 59.176, 59.1649, 59.1647, 59.1594, 
    59.1569, 59.1613, 59.1622, 59.1679, 59.1745, 59.1798, 59.2189, 59.2256, 
    59.2264, 59.2326, 59.2319, 59.2322, 59.2302, 59.2257, 59.2264, 59.2223, 
    59.2301, 59.222, 59.2184, 59.2181, 59.2223, 59.2269, 59.2219, 59.221, 
    59.2257, 59.224, 59.2269, 59.2238, 59.2252, 59.2267, 59.2254, 59.2276, 
    59.2256, 59.2253, 59.2202, 59.2267, 59.226, 59.2221, 59.2169, 59.2163, 
    59.2261, 59.2256, 59.2257, 59.213, 59.208, 59.204, 59.2072, 59.2054, 
    59.2065, 59.206, 59.2023, 59.2025, 59.207, 59.2065, 59.2066, 59.1719, 
    59.1523, 59.1485, 59.1016, 59.101, 59.0923, 59.1003, 59.1004, 59.1011, 
    59.0801, 59.0942, 59.0939, 59.0853, 59.0913, 59.0926, 59.092, 59.0989, 
    59.096, 59.0979, 59.0967, 59.0954, 59.095, 59.0922, 59.0864, 59.0882, 
    59.0991, 59.1979, 58.9858, 59.1626, 59.1612, 59.1546, 59.1445, 59.1429, 
    59.1315, 59.1205, 59.1421, 59.1221, 59.1317, 59.1315, 59.1315, 59.1322, 
    59.1315, 59.1306, 59.1249, 59.1285, 59.1296, 59.129, 59.1318, 59.1304, 
    59.1274, 59.1269, 59.1286, 59.1182, 59.0948, 59.0977, 59.1191, 59.1229, 
    59.1348, 59.1337, 59.1463, 59.1414, 59.1781, 59.1747, 59.1885, 59.1925, 
    59.2001, 59.1984, 59.1745, 59.1592, 59.182, 59.1908, 59.1773, 59.2116, 
    59.2116, 59.2051, 59.2079, 59.2059, 59.2119, 59.2069, 59.2062, 59.2071, 
    59.2034, 59.206, 59.204, 59.2054, 59.2078, 59.2043, 59.198, 59.2001, 
    59.1974, 59.192, 59.1947, 59.1954, 59.1843, 59.1657, 59.229, 59.2137, 
    59.2099, 59.2099, 59.2097, 59.1871, 59.1751, 59.1686, 59.1838, 59.1768, 
    59.1882, 59.1633, 59.1685, 59.1856, 59.1988, 59.1887, 59.2013, 59.1902, 
    59.1897, 59.2138, 59.2133, 59.2024, 59.2099, 59.1922, 59.1945, 59.1951, 
    59.1924, 59.1964, 59.192, 59.1918, 59.1901, 59.1926, 59.1943, 59.1951, 
    59.195, 59.1964, 59.1966, 59.1911, 59.1938, 59.2001, 59.1869, 59.1812, 
    59.1956, 59.218, 59.1948, 59.2337, 59.2427, 59.2302, 59.1983, 59.1969, 
    59.1929, 59.1909, 59.1911, 59.1955, 59.1889, 59.1958, 59.1947, 59.1956, 
    59.1946, 59.1829, 59.1911, 59.1914, 59.1922, 59.1948, 59.1683, 59.1708, 
    59.1727, 59.1427, 59.1423, 59.1358, 59.1413, 59.1235, 59.1207, 59.1196, 
    59.1193, 59.1313, 59.1188, 59.1178, 59.1324, 59.1335, 59.137, 59.1331, 
    59.1364, 59.1362, 59.1333, 59.1312, 59.1465, 59.1505, 59.1628, 59.1623, 
    59.1538, 59.1276, 59.1167, 59.0935, 59.0952, 59.0685, 59.0954, 59.1, 
    59.0973, 59.0884, 59.128, 59.1246, 59.1272, 59.1242, 59.1217, 59.1256, 
    59.1229, 59.1107, 59.1138, 59.1109, 59.0992, 59.0973, 59.096, 59.0934, 
    59.0952, 59.0955, 59.0946, 59.0951, 59.0952, 59.1162, 59.0885, 59.0796, 
    59.1042, 59.1057, 59.1074, 59.0991, 59.0991, 59.1029, 59.1331, 59.1354, 
    59.1308, 59.1384, 59.1312, 59.1475, 59.1521, 59.1536, 59.1731, 59.1663, 
    59.1723, 59.1706, 59.1957, 59.1955, 59.1914, 59.191, 59.1842, 59.2214, 
    59.2179, 59.2118, 59.2593, 59.2152, 59.2037, 59.2028, 59.2335, 59.1899, 
    59.2149, 59.2267, 59.2545, 59.2533, 59.2549, 59.2486, 59.2553, 59.2416, 
    59.2377, 59.2242, 59.1972, 59.2073, 59.2064, 59.1924, 59.1932, 59.1698, 
    59.1933, 59.1873, 59.193, 59.1708, 59.1956, 59.1912, 59.2215, 59.2276, 
    59.2233, 59.2337, 59.2311, 59.2311, 59.232, 59.2403, 59.2438, 59.2415, 
    59.2263, 59.2428, 59.2426, 59.2441, 59.2455, 59.2321, 59.2405, 59.2406, 
    59.2259, 59.2429, 59.2433, 59.241, 59.2436, 59.2412, 59.2578, 59.2408, 
    59.2401, 59.2399, 59.2415, 59.2415, 59.2315, 59.2315, 59.2327, 59.2387, 
    59.2383, 59.2484, 59.2479, 59.237, 59.2378, 59.2225, 59.2388, 59.2447, 
    59.237, 59.2377, 59.24, 59.2325, 59.2385, 59.2367, 59.2402, 59.2376, 
    59.2337, 59.2408, 59.2335, 59.2354, 59.236, 59.2355, 59.236, 59.2359, 
    59.2377, 59.2373, 59.239, 59.2433, 59.2415, 59.2415, 59.244, 59.2426, 
    59.247, 59.2439, 59.2472, 59.2492, 59.2493, 59.2483, 59.2509, 59.2493, 
    59.2424, 59.2426, 59.2424, 59.2405, 59.2453, 59.2316, 59.2341, 59.246, 
    59.2421, 59.2454, 59.2463, 59.2408, 59.2425, 59.2478, 59.2408, 59.2474, 
    59.2406, 59.2407, 59.2367, 59.2359, 59.2355, 59.2439, 59.244, 59.2437, 
    59.2441, 59.241, 59.2422, 59.2405, 59.2476, 59.2439, 59.2507, 59.2466, 
    59.2431, 59.2448, 59.2454, 59.234, 59.2202, 59.236, 59.2332, 59.2216, 
    59.2265, 59.2455, 59.2428, 59.2411, 59.1962, 59.2559, 59.2419, 59.2385, 
    59.2393, 59.2388, 59.2427, 59.2425, 59.2398, 59.2382, 59.2379, 59.2364, 
    59.2388, 59.2421, 59.2362, 59.2363, 59.235, 59.2313, 59.2333, 59.2314, 
    59.2271, 59.2378, 59.2369, 59.2366, 59.2181, 59.2436, 59.2442, 59.2442, 
    59.2418, 59.2404, 59.2438, 59.2396, 59.2347, 59.2268, 59.2267, 59.2278, 
    59.2235, 59.2248, 59.2252, 59.2408, 59.2402, 59.2294, 59.2343, 59.2326, 
    59.24, 59.2367, 59.2376, 59.237, 59.2378, 59.2351, 59.2309, 59.2139, 
    59.1996, 59.1793, 59.2012, 59.2044, 59.192, 59.2033, 59.209, 59.2033, 
    59.2083, 59.2079, 59.2586, 59.2493, 59.2261, 59.226, 59.2227, 59.2425, 
    59.2365, 59.2453, 59.253, 59.2379, 59.2366, 59.2405, 59.2448, 59.2391, 
    59.2376, 59.2376, 59.2301, 59.2275, 59.2294, 59.1932, 59.2153, 59.228, 
    59.2282, 59.2289, 59.232, 59.2384, 59.2508, 59.239, 59.2472, 59.2424, 
    59.2415, 59.2357, 59.2421, 59.2466, 59.2518, 59.2517, 59.2503, 59.2521, 
    59.2503, 59.2319, 59.2683, 59.2732, 59.2533, 59.2585, 59.2543, 59.2528, 
    59.2466, 59.2356, 59.2464, 59.2387, 59.2446, 59.2361, 59.2416, 59.2468, 
    59.2397, 59.239, 59.2387, 59.246, 59.2536, 59.2418, 59.2401, 59.2351, 
    59.2331, 59.2418, 59.2589, 59.2835, 59.2795, 59.2722, 59.1504, 59.1467, 
    59.1393, 59.1377, 59.1338, 59.1367, 59.137, 59.1126, 59.1153, 59.1128, 
    59.1001, 59.0992, 59.0978, 59.0919, 59.1029, 59.1002, 59.0936, 59.0951, 
    59.0952, 59.0827, 59.0953, 59.0977, 59.1304, 59.1367, 59.1277, 59.0928, 
    59.0931, 59.0754, 59.0948, 59.0951, 59.095, 59.0997, 59.0959, 59.0954, 
    59.0931, 59.0928, 59.0714, 59.0849, 59.0804, 59.1006, 59.0861, 59.0925, 
    59.0878, 59.1124, 59.1138, 59.1301, 59.1236, 59.1228, 59.1412, 59.1194, 
    59.1545, 59.1202, 59.163, 59.153, 59.1628, 59.1752, 59.1844, 59.1932, 
    59.1938, 59.1958, 59.2005, 59.2051, 59.1532, 59.16, 59.1557, 59.1667, 
    59.2476, 59.2014, 59.196, 59.1656, 59.2319, 59.2401, 59.2655, 59.3085, 
    59.2731, 59.217, 59.2285, 59.2286, 59.2324, 59.2383, 59.2289, 59.231, 
    59.2385, 59.2328, 59.2129, 59.2146, 59.1931, 59.2147, 59.2206, 59.236, 
    59.2395, 59.2415, 59.2531, 59.242, 59.2495, 59.2432, 59.236, 59.2165, 
    59.2234, 59.2173, 59.1997, 59.2243, 59.2001, 59.223, 59.2233, 59.1954, 
    59.1557, 59.1724, 59.1772, 59.1817, 59.1964, 59.1963, 59.1704, 59.1863, 
    59.1859, 59.1859, 59.1856, 59.1858, 59.2022, 59.1868, 59.1956, 59.1965, 
    59.1853, 59.1866, 59.1862, 59.2182, 59.2201, 59.2239, 59.2237, 59.2253, 
    59.2261, 59.2275, 59.2266, 59.2266, 59.2275, 59.2273, 59.226, 59.2257, 
    59.181, 59.2232, 59.1861, 59.193, 59.2046, 59.2209, 59.2087, 59.209, 
    59.2086, 59.2138, 59.2067, 59.1938, 59.1954, 59.1925, 59.2139, 59.2112, 
    59.1816, 59.1947, 59.1729, 59.163, 59.1632, 59.1643, 59.1515, 59.1702, 
    59.1725, 59.1747, 59.1739, 59.1763, 59.1769, 59.1934, 59.1768, 59.1764, 
    59.1762, 59.1765, 59.2088, 59.2195, 59.2228, 59.2299, 59.225, 59.2514, 
    59.2471, 59.2487, 59.244, 59.2405, 59.2399, 59.2275, 59.2234, 59.2235, 
    59.2233, 59.2149, 59.2018, 59.1963, 59.1959, 59.1931, 59.1943, 59.1937, 
    59.1936, 59.1883, 59.1933, 59.193, 59.1799, 59.19, 59.19, 59.1864, 
    59.1898, 59.1937, 59.1945, 59.1941, 59.1897, 59.2006, 59.1972, 59.2023, 
    59.1916, 59.1783, 59.1835, 59.1962, 59.2161, 59.188, 59.1887, 59.222, 
    59.2157, 59.2077, 59.2171, 59.2105, 59.2174, 59.2023, 59.196, 59.2013, 
    59.2065, 59.175, 59.1592, 59.1652, 59.1651, 59.1568, 59.1335, 59.1275, 
    59.1056, 59.0935, 59.0909, 59.0957, 59.0954, 59.0872, 59.097, 59.0949, 
    59.0952, 59.0937, 59.0458, 59.0936, 59.0804, 59.095, 59.0908, 59.0893, 
    59.0905, 59.0948, 59.0943, 59.094, 59.0961, 59.0964, 59.0955, 59.0955, 
    59.0821, 59.0877, 59.0943, 59.0944, 59.095, 59.0923, 59.0938, 59.095, 
    59.0944, 59.1008, 59.1111, 59.1196, 59.1191, 59.1219, 59.1595, 59.1632, 
    59.1632, 59.1629, 59.1811, 59.1762, 59.1796, 59.1776, 59.199, 59.1959, 
    59.1702, 59.1776, 59.1786, 59.159, 59.1765, 59.0775, 59.0706, 59.0701, 
    59.178, 59.1746, 59.0923, 59.0927, 59.0915, 59.0972, 59.1138, 59.1009, 
    59.1313, 59.1295, 59.1122, 59.1802, 59.1856, 59.194, 59.1934, 59.1968, 
    59.191, 59.1912, 59.1931, 59.1939, 59.2039, 59.2008, 59.1933, 59.1933, 
    59.1926, 59.1988, 59.192, 59.1931, 59.1957, 59.1938, 59.1938, 59.1954, 
    59.1932, 59.2009, 59.2029, 59.2068, 59.2368, 59.221, 59.2223, 59.2209, 
    59.2234, 59.1948, 59.2223, 59.223, 59.186, 59.258, 59.2495, 59.2496, 
    59.2504, 59.2505, 59.2332, 59.2687, 59.2554, 59.2568, 59.26, 59.2483, 
    59.2614, 59.2677, 59.2231, 59.2705, 59.2186, 59.2115, 59.2523, 59.2017, 
    59.1943, 59.1912, 59.1974, 59.1968, 59.1943, 59.1746, 59.1712, 59.1592, 
    59.1489, 59.1619, 59.1417, 59.1797, 59.1788, 59.1773, 59.2276, 59.2108, 
    59.2314, 59.2105, 59.2043, 59.2013, 59.2104, 59.2124, 59.2104, 59.2092, 
    59.2108, 59.2093, 59.2089, 59.2109, 59.2138, 59.2187, 59.2209, 59.2209, 
    59.2179, 59.2118, 59.2101, 59.2191, 59.2228, 59.2148, 59.209, 59.2106, 
    59.2132, 59.2099, 59.2049, 59.2104, 59.2121, 59.2237, 59.2231, 59.2242, 
    59.2222, 59.2215, 59.2348, 59.2095, 59.2104, 59.1985, 59.1911, 59.1965, 
    59.1953, 59.2001, 59.2044, 59.2104, 59.2102, 59.1843, 59.1953, 59.1946, 
    59.1953, 59.1976, 59.1883, 59.1955, 59.1951, 59.1969, 59.2004, 59.1936, 
    59.1909, 59.1935, 59.2004, 59.2004, 59.1967, 59.1992, 59.1926, 59.182, 
    59.2002, 59.1995, 59.1963, 59.1957, 59.1962, 59.1959, 59.1965, 59.1961, 
    59.1983, 59.1959, 59.1941, 59.1957, 59.1976, 59.2007, 59.1919, 59.2006, 
    59.1964, 59.1957, 59.1948, 59.1954, 59.2001, 59.1963, 59.1936, 59.195, 
    59.1953, 59.1947, 59.198, 59.1962, 59.1978, 59.1978, 59.1958, 59.186, 
    59.1932, 59.1962, 59.1962, 59.1979, 59.1986, 59.1958, 59.1837, 59.2121, 
    59.2057, 59.205, 59.2247, 59.204, 59.2027, 59.1859, 59.1852, 59.1858, 
    59.1808, 59.1885, 59.1918, 59.1926, 59.1925, 59.1935, 59.1947, 59.1923, 
    59.1904, 59.1738, 59.1693, 59.1639, 59.1619, 59.1459, 59.1441, 59.1501, 
    59.1526, 59.1494, 59.1395, 59.0892, 59.0946, 59.0957, 59.0196, 59.085, 
    59.075, 59.0942, 59.098, 59.0936, 59.0886, 59.095, 59.0932, 59.0902, 
    59.0971, 59.097, 59.0895, 59.0949, 59.0943, 59.095, 59.0966, 59.0942, 
    59.0933, 59.1045, 59.1036, 59.12, 59.2328, 59.1968, 59.2059, 59.2044, 
    59.206, 59.2165, 59.2122, 59.2038, 59.1968, 59.1242, 59.1017, 59.0967, 
    59.0977, 59.0938, 59.0945, 59.092, 59.0919, 59.0815, 59.0945, 59.0805, 
    59.0889, 59.0926, 59.0953, 59.0962, 59.095, 59.0925, 59.0975, 59.099, 
    59.0877, 59.0857, 59.0903, 59.0914, 59.0911, 59.0901, 59.0895, 59.0919, 
    59.0951, 59.0906, 59.0906, 59.0906, 59.1005, 59.1136, 59.1624, 59.1595, 
    59.1944, 59.1978, 59.0804, 59.1419, 59.1916, 59.1839, 59.1527, 59.1808, 
    59.1724, 59.1402, 59.1545, 59.1565, 59.1941, 59.1918, 59.2044, 59.2005, 
    59.2022, 59.1942, 59.1989, 59.1998, 59.1942, 59.203, 59.194, 59.1961, 
    59.1961, 59.1981, 59.1985, 59.1956, 59.1948, 59.2013, 59.1967, 59.1933, 
    59.2058, 59.2224, 59.1937, 59.1962, 59.1966, 59.1963, 59.1965, 59.1965, 
    59.2923, 59.2092, 59.2101, 59.2213, 59.2131, 59.2125, 59.2169, 59.2117, 
    59.2103, 59.2229, 59.1979, 59.2097, 59.2235, 59.2239, 59.2107, 59.2117, 
    59.209, 59.2114, 59.2091, 59.2118, 59.2111, 59.2128, 59.1943, 59.2084, 
    59.2112, 59.2073, 59.2076, 59.2069, 59.2077, 59.2087, 59.2082, 59.2127, 
    59.2223, 59.2227, 59.2219, 59.2214, 59.2218, 59.2245, 59.2528, 59.2255, 
    59.2481, 59.226, 59.2103, 59.2453, 59.2071, 59.1911, 59.1902, 59.1821, 
    59.1869, 59.1773, 59.1812, 59.181, 59.1807, 59.181, 59.1808, 59.1848, 
    59.196, 59.1959, 59.1959, 59.1961, 59.1961, 59.1966, 59.1962, 59.1875, 
    59.1841, 59.1956, 59.1957, 59.1972, 59.1976, 59.1965, 59.2195, 59.2206, 
    59.2227, 59.2117, 59.2115, 59.2123, 59.2101, 59.2166, 59.2096, 59.2235, 
    59.2091, 59.211, 59.2118, 59.2068, 59.1859, 59.1976, 59.1982, 59.1849, 
    59.2041, 59.2369, 59.1893, 59.1793, 59.1721, 59.1643, 59.2606, 59.0911, 
    59.0925, 59.0917, 59.0945, 59.0951, 59.0945, 59.0947, 59.0895, 59.0938, 
    59.0961, 59.0963, 59.0958, 59.0964, 59.0967, 59.0942, 59.0944, 59.0957, 
    59.0948, 59.0956, 59.0918, 59.0939, 59.0863, 59.2042, 59.2049, 59.2053, 
    59.2061, 59.2064, 59.2117, 59.2043, 59.203, 59.2022, 59.199, 59.2006, 
    59.2008, 59.2062, 59.2118, 59.1948, 59.2086, 59.2078, 59.2066, 59.2131, 
    59.2247, 59.2197, 59.2202, 59.2242, 59.2238, 59.2206, 59.2055, 59.2025, 
    59.2018, 59.2029, 59.184, 59.1857, 59.1863, 59.1858, 59.1907, 59.1928, 
    59.1921, 59.1982, 59.1982, 59.1874, 59.1882, 59.1475, 59.1922, 59.161, 
    59.1811, 59.195, 59.1922, 59.1968, 59.1984, 59.198, 59.1956, 59.198, 
    59.2022, 59.1957, 59.2002, 59.2048, 59.2126, 59.1973, 59.1964, 59.2086, 
    59.2046, 59.2089, 59.2017, 59.2189, 59.1931, 59.1885, 59.1924, 59.1928, 
    59.19, 59.1859, 59.1892, 59.1756, 59.1814, 59.1928, 59.2001, 59.2, 
    59.1996, 59.1294, 59.2021, 59.201, 59.2003, 59.1984, 59.1984, 59.1987, 
    59.1982, 59.1985, 59.2024, 59.196, 59.1958, 59.1982, 59.1989, 59.199, 
    59.1983, 59.1924, 59.1883, 59.1848, 59.1794, 59.1698, 59.1822, 59.1847, 
    59.1876, 59.1866, 59.1848, 59.1848, 59.1894, 59.2012, 59.2015, 59.2015, 
    59.2023, 59.1976, 59.1703, 59.2057, 59.1713, 59.1737, 59.1779, 59.1726, 
    59.1748, 59.1753, 59.1792, 59.171, 59.2003, 59.1755, 59.1712, 59.1778, 
    59.1823, 59.1798, 59.1876, 59.1963, 59.2049, 59.1528, 59.2193, 59.2224, 
    59.2243, 59.2328, 59.2229, 59.2196, 59.2201, 59.2201, 59.2191, 59.2111, 
    59.2205, 59.2164, 59.2091, 59.1969, 59.1857, 59.2136, 59.177, 59.1738, 
    59.1618, 59.1697, 59.1626, 59.1461, 59.1413, 59.0998, 59.1341, 59.1322, 
    59.1252, 59.1238, 59.1138, 59.1211, 59.1226, 59.0952, 59.0934, 59.1208, 
    59.1221, 59.1969, 59.2227, 59.2214, 59.1688, 59.1705, 59.1673, 59.1718, 
    59.1608, 59.176, 59.1662, 59.1721, 59.182, 59.1562, 59.1759, 59.1671, 
    59.1621, 59.1627, 59.1791, 59.1775, 59.1796, 59.1877, 59.1851, 59.196, 
    59.1866, 59.188, 59.222, 59.1734, 59.192, 59.1466, 59.1564, 59.1601, 
    59.1651, 59.1734, 59.1751, 59.1625, 59.1601, 59.1583, 59.2171, 59.2137, 
    59.2131, 59.2157, 59.22, 59.2355, 59.2178, 59.2284, 59.2279, 59.2296, 
    59.2286, 59.2294, 59.2157, 59.2164, 59.2097, 59.2078, 59.2004, 59.2124, 
    59.2123, 59.2112, 59.2115, 59.2121, 59.2116, 59.2079, 59.2104, 59.2092, 
    59.1939, 59.1868, 59.194, 59.2129, 59.2776, 59.2736, 59.2179, 59.2214, 
    59.2113, 59.2208, 59.2285, 59.2133, 59.2144, 59.2184, 59.2204, 59.2333, 
    59.2245, 59.2252, 59.2277, 59.1925, 59.1933, 59.195, 59.2089, 59.199, 
    59.1809, 59.1811, 59.1907, 59.1902, 59.191, 59.1877, 59.1909, 59.1908, 
    59.2046, 59.2206, 59.21, 59.2112, 59.2156, 59.2243, 59.2224, 59.2172, 
    59.2273, 59.2091, 59.1925, 59.1819, 59.1836, 59.1839, 59.2027, 59.125, 
    59.125, 59.1303, 59.1074, 59.0948, 59.0956, 59.0942, 59.0849, 59.1054, 
    59.0934, 59.0949, 59.0993, 59.0932, 59.0986, 59.0967, 59.0955, 59.0951, 
    59.0942, 59.0937, 59.0947, 59.0955, 59.0993, 59.0983, 59.0965, 59.1005, 
    59.1057, 59.18, 59.0912, 59.1759, 59.1758, 59.1504, 59.1445, 59.1503, 
    59.1582, 59.1436, 59.1368, 59.1003, 59.1228, 59.123, 59.1169, 59.1004, 
    59.1035, 59.104, 59.1029, 59.0738, 59.1061, 59.1119, 59.1077, 59.1021, 
    59.0978, 59.0851, 59.102, 59.1023, 59.0968, 59.0969, 59.1, 59.0979, 
    59.0989, 59.0941, 59.0937, 59.0964, 59.0981, 59.0972, 59.0992, 59.1104, 
    59.1173, 59.1448, 59.1515, 59.1712, 59.1825, 59.1882, 59.1806, 59.1639, 
    59.1669, 59.1779, 59.1696, 59.1589, 59.1559, 59.1636, 59.1786, 59.1911, 
    59.0777, 59.1771, 59.2037, 59.2033, 59.1954, 59.2009, 59.1961, 59.1998, 
    59.1973, 59.1997, 59.2001, 59.2063, 59.2039, 59.2051, 59.2073, 59.219, 
    59.2446, 59.2421, 59.2567, 59.2244, 59.1795, 59.1825, 59.1694, 59.2095, 
    59.1937, 59.152, 59.1963, 59.1922, 59.2076, 59.2054, 59.2006, 59.1983, 
    59.1971, 59.1929, 59.1933, 59.193, 59.1949, 59.1963, 59.1942, 59.1975, 
    59.1984, 59.1983, 59.1968, 59.1956, 59.1954, 59.1957, 59.1959, 59.1938, 
    59.196, 59.1959, 59.1906, 59.1922, 59.1986, 59.2002, 59.1992, 59.1965, 
    59.1957, 59.1958, 59.1955, 59.1954, 59.196, 59.1957, 59.1953, 59.1957, 
    59.1959, 59.1961, 59.1977, 59.1962, 59.2006, 59.2001, 59.2061, 59.2061, 
    59.212, 59.2128, 59.2142, 59.2151, 59.2137, 59.2124, 59.2102, 59.2124, 
    59.2101, 59.2226, 59.2197, 59.2275, 59.2247, 59.2174, 59.2217, 59.216, 
    59.1926, 59.2106, 59.2018, 59.2084, 59.2086, 59.2077, 59.1782, 59.2012, 
    59.2021, 59.1964, 59.2228, 59.2168, 59.2285, 59.2275, 59.226, 59.2344, 
    59.2304, 59.2263, 59.2262, 59.2264, 59.2252, 59.2135, 59.2177, 59.2193, 
    59.205, 59.2022, 59.1974, 59.1874, 59.2073, 59.1857, 59.1876, 59.191, 
    59.1662, 59.1743, 59.166, 59.1608, 59.1195, 59.1328, 59.1096, 59.0938, 
    59.0888, 59.0951, 59.0951, 59.0874, 59.0949, 58.7985, 59.0929, 59.0973, 
    59.0965, 59.0947, 59.0925, 59.0964, 59.0963, 59.0956, 59.0929, 59.0929, 
    59.0943, 59.0953, 59.0966, 59.0969, 59.0979, 59.1103, 59.1235, 59.1245, 
    59.1284, 59.1463, 59.1312, 59.1293, 59.1547, 59.1647, 59.1638, 59.1718, 
    59.1716, 59.1744, 59.176, 59.198, 59.1925, 59.1946, 59.2012, 59.1952, 
    59.1992, 59.2066, 59.1945, 59.2092, 59.1952, 59.1857, 59.1899, 59.1923, 
    59.1907, 59.1944, 59.1835, 59.1812, 59.1645, 59.1646, 59.1627, 59.1633, 
    59.2096, 59.1837, 59.1894, 59.1887, 59.1834, 59.1817, 59.1822, 59.1874, 
    59.18, 59.1749, 59.1748, 59.1716, 59.1691, 59.1701, 59.1703, 59.1756, 
    59.1888, 59.1812, 59.2029, 59.1964, 59.2028, 59.2051, 59.1842, 59.2086, 
    59.1963, 59.1876, 59.1799, 59.1781, 59.189, 59.197, 59.203, 59.1687, 
    59.1942, 59.1917, 59.1833, 59.1812, 59.2065, 59.1562, 59.1694, 59.2066, 
    59.2066, 59.2026, 59.2279, 59.228, 59.228, 59.2275, 59.2275, 59.229, 
    59.2283, 59.2284, 59.2272, 59.2265, 59.2234, 59.2268, 59.2377, 59.2366, 
    59.2318, 59.2318, 59.2305, 59.2305, 59.188, 59.2009, 59.2072, 59.2043, 
    59.1946, 59.1874, 59.131, 59.1341, 59.1303, 59.1956, 59.2012, 59.1974, 
    59.2004, 59.2001, 59.2, 59.2011, 59.2062, 59.2024, 59.1954, 59.2162, 
    59.2227, 59.1768, 59.2144, 59.2337, 59.2224, 59.2331, 59.2152, 59.2091, 
    59.2092, 59.2092, 59.3466, 59.18, 59.181, 59.1768, 59.1874, 59.1875, 
    59.1852, 59.1849, 59.1852, 59.192, 59.1952, 59.2019, 59.1803, 59.1832, 
    59.1814, 59.1857, 59.1812, 59.1814, 59.1819, 59.1744, 59.1888, 59.1762, 
    59.1774, 59.168, 59.1747, 59.0922, 59.1082, 59.118, 59.1276, 59.1163, 
    59.1125, 59.1618, 59.1653, 59.166, 59.1857, 59.1853, 59.1853, 59.195, 
    59.1956, 59.199, 59.2001, 59.1999, 59.2, 59.198, 59.2033, 59.1804, 
    59.1841, 59.1964, 59.2034, 59.2094, 59.2097, 59.2096, 59.2097, 59.2307, 
    59.2091, 59.2052, 59.2071, 59.2069, 59.2064, 59.206, 59.2057, 59.1944, 
    59.1709, 59.2022, 59.2202, 59.2205, 59.2117, 59.199, 59.1966, 59.1934, 
    59.1947, 59.1985, 59.1986, 59.1974, 59.1964, 59.1972, 59.1954, 59.1995, 
    59.1993, 59.1969, 59.1983, 59.1975, 59.2007, 59.1937, 59.1964, 59.1982, 
    59.1959, 59.1951, 59.1979, 59.1966, 59.1979, 59.1931, 59.1927, 59.1996, 
    59.1996, 59.198, 59.1891, 59.1936, 59.1754, 59.1773, 59.1915, 59.1996, 
    59.1993, 59.2003, 59.1996, 59.2004, 59.1645, 59.1978, 59.1786, 59.1765, 
    59.1772, 59.1749, 59.1762, 59.1893, 59.2057, 59.2057, 59.1943, 59.1928, 
    59.1943, 59.1799, 59.1992, 59.1982, 59.1968, 59.1972, 59.1987, 59.1987, 
    59.2031, 59.1957, 59.1969, 59.1983, 59.2037, 59.1978, 59.1994, 59.1997, 
    59.1996, 59.1991, 59.2093, 59.1998, 59.1814, 59.1795, 59.214, 59.2383, 
    59.2109, 59.2195, 59.2143, 59.2195, 59.2155, 59.2157, 59.2205, 59.2218, 
    59.2206, 59.2203, 59.2277, 59.2276, 59.2196, 59.2182, 59.2199, 59.2168, 
    59.2119, 59.2128, 59.219, 59.219, 59.219, 59.2186, 59.2185, 59.2223, 
    59.2188, 59.2184, 59.1976, 59.1849, 59.1866, 59.1823, 59.1248, 59.1144, 
    59.099, 59.1093, 59.1258, 59.1213, 59.1259, 59.1279, 59.1294, 59.1303, 
    59.1285, 59.1283, 59.1283, 59.1288, 59.1218, 59.1105, 59.1249, 59.1027, 
    59.1149, 59.0975, 59.0858, 59.0953, 59.0962, 59.0951, 59.0954, 59.0952, 
    59.096, 59.0927, 59.0973, 59.0978, 59.0979, 59.1111, 58.9208, 59.1182, 
    59.0758, 59.1623, 59.1631, 59.159, 59.1957, 59.1923, 59.2108, 59.217, 
    59.2527, 59.2243, 59.2265, 59.2367, 59.2384, 59.225, 59.2294, 59.2205, 
    59.2187, 59.2269, 59.2202, 59.2189, 59.2186, 59.2148, 59.2203, 59.2193, 
    59.2181, 59.2236, 59.2186, 59.2188, 59.219, 59.2199, 59.2189, 59.2283, 
    59.2278, 59.2198, 59.2186, 59.2123, 59.2147, 59.2044, 59.1985, 59.1969, 
    59.1955, 59.1995, 59.1988, 59.2028, 59.1937, 59.1966, 59.1987, 59.1931, 
    59.1989, 59.1995, 59.1976, 59.1989, 59.196, 59.1921, 59.1956, 59.1919, 
    59.198, 59.1987, 59.1905, 59.2047, 59.2045, 59.1844, 59.1706, 59.1669, 
    59.2103, 59.2015, 59.2157, 59.2215, 59.2163, 59.2227, 59.203, 59.1872, 
    59.1994, 59.1995, 59.2002, 59.2015, 59.1857, 59.1855, 59.1781, 59.1846, 
    59.1863, 59.1995, 59.1994, 59.1785, 59.1681, 59.1662, 59.1665, 59.1884, 
    59.165, 59.2229, 59.233, 59.2419, 59.2503, 59.1928, 59.1936, 59.253, 
    59.2053, 59.2142, 59.2185, 59.2226, 59.2214, 59.2031, 59.2123, 59.2115, 
    59.2124, 59.2117, 59.1945, 59.2173, 59.2336, 59.2242, 59.2029, 59.2128, 
    59.2175, 59.2098, 59.2118, 59.2098, 59.2145, 59.2045, 59.1966, 59.1931, 
    59.2128, 59.2078, 59.2167, 59.212, 59.2122, 59.2084, 59.2006, 59.2064, 
    59.1937, 59.1771, 59.1683, 59.1723, 59.1808, 59.1789, 59.1869, 59.1989, 
    59.1829, 59.1811, 59.1812, 59.1953, 59.2061, 59.1913, 59.1961, 59.1937, 
    59.2122, 59.216, 59.2165, 59.2079, 59.1869, 59.2011, 59.2092, 59.1961, 
    59.215, 59.1803, 59.2108, 59.2085, 59.1875, 59.2122, 59.2147, 59.184, 
    59.1818, 59.1881, 59.2026, 59.2019, 59.2099, 59.2187, 59.2046, 59.2051, 
    59.1992, 59.1984, 59.1959, 59.1947, 59.1974, 59.1951, 59.2047, 59.2003, 
    59.2005, 59.1958, 59.2153, 59.1957, 59.2071, 59.2024, 59.203, 59.2016, 
    59.2016, 59.2129, 59.2146, 59.2107, 59.2103, 59.2152, 59.2157, 59.2204, 
    59.192, 59.2358, 59.2276, 59.1797, 59.1817, 59.1777, 59.1798, 59.1651, 
    59.1644, 59.1963, 59.1646, 59.18, 59.183, 59.21, 59.1928, 59.1857, 
    59.1978, 59.1973, 59.1976, 59.1954, 59.1967, 59.1854, 59.1881, 59.1884, 
    59.1951, 59.1842, 59.1747, 59.1797, 59.1783, 59.1783, 59.1838, 59.1863, 
    59.1854, 59.1863, 59.2017, 59.1944, 59.1907, 59.1867, 59.1695, 59.1889, 
    59.1344, 59.1416, 59.1728, 59.1623, 59.1602, 59.1926, 59.1861, 59.1926, 
    59.1874, 59.1723, 59.1386, 59.1354, 59.1284, 59.1188, 59.1165, 59.1996, 
    59.1108, 59.1053, 59.1034, 59.0846, 59.0938, 59.0985, 59.0946, 59.0993, 
    59.0958, 59.0953, 59.0906, 59.0941, 59.0936, 59.0936, 59.0952, 59.0966, 
    59.0963, 59.0944, 59.0937, 59.0943, 59.0955, 59.0992, 59.0944, 59.0946, 
    59.095, 59.0953, 59.0941, 59.0904, 59.0089, 59.0225, 59.2062, 59.2072, 
    59.2077, 59.2205, 59.2034, 59.2047, 59.2035, 59.2042, 59.2066, 59.2063, 
    59.2102, 59.2094, 59.2133, 59.2017, 59.2021, 59.1955, 59.1977, 59.1848, 
    59.2061, 59.2058, 59.2042, 59.2248, 59.2269, 59.228, 59.2198, 59.1803, 
    59.2151, 59.1614, 59.1767, 59.1854, 59.1768, 59.1934, 59.1952, 59.228, 
    59.2272, 59.212, 59.2089, 59.2195, 59.2256, 59.2194, 59.2228, 59.2207, 
    59.2165, 59.2173, 59.2187, 59.219, 59.2116, 59.2153, 59.2205, 59.2865, 
    59.2231, 59.2236, 59.2235, 59.3443, 59.2235, 59.2189, 59.2183, 59.2196, 
    59.2139, 59.2039, 59.1843, 59.1774, 59.1706, 59.1815, 59.1742, 59.1779, 
    59.1764, 59.2137, 59.3227, 59.3137, 59.1917, 59.1899, 59.2044, 59.1925, 
    59.2135, 59.2167, 59.2119, 59.1996, 59.2081, 59.2098, 59.2054, 59.2126, 
    59.21, 59.2125, 59.2125, 59.2128, 59.2118, 59.2126, 59.2142, 59.2183, 
    59.222, 59.2211, 59.2254, 59.2208, 59.2507, 59.2541, 59.2344, 59.2158, 
    59.2105, 59.1929, 59.1967, 59.1447, 59.1811, 59.186, 59.1788, 59.1646, 
    59.1484, 59.1794, 59.1794, 59.1832, 59.1706, 59.1683, 59.1909, 59.1736, 
    59.1819, 59.1795, 59.1679, 59.1794, 59.1672, 59.1695, 59.198, 59.1974, 
    59.1992, 59.1983, 59.1816, 59.2023, 59.1995, 59.1995, 59.199, 59.1963, 
    59.1666, 59.1729, 59.2615, 59.1883, 59.1901, 59.1717, 59.1645, 59.1594, 
    59.1548, 59.105, 59.1, 59.0926, 59.0947, 59.0943, 59.0901, 59.094, 
    59.0938, 59.0941, 59.0901, 59.0921, 59.0955, 59.0942, 59.0945, 59.0968, 
    59.0939, 59.0923, 59.0969, 59.0924, 59.0931, 59.0955, 59.0966, 59.092, 
    59.0701, 59.1101, 59.1296, 59.1475, 59.1654, 59.1598, 59.174, 59.1751, 
    59.185, 59.1861, 59.1836, 59.1844, 59.1786, 59.1828, 59.1839, 59.1813, 
    59.1805, 59.1816, 59.1874, 59.1856, 59.188, 59.1899, 59.192, 59.2019, 
    59.2033, 59.1623, 59.1687, 59.1864, 59.1785, 59.1784, 59.1854, 59.1882, 
    59.1864, 59.1771, 59.1743, 59.182, 59.1793, 59.1828, 59.179, 59.1926, 
    59.1977, 59.1959, 59.195, 59.1978, 59.1938, 59.2119, 59.1912, 59.1969, 
    59.1872, 59.2, 59.1958, 59.1969, 59.1973, 59.1912, 59.1954, 59.1893, 
    59.1701, 59.159, 59.161, 59.1661, 59.1728, 59.165, 59.1595, 59.1806, 
    59.1587, 59.1542, 59.1613, 59.1643, 59.1698, 59.1682, 59.1861, 59.1871, 
    59.1863, 59.173, 59.1738, 59.1779, 59.1829, 59.1827, 59.1804, 59.1857, 
    59.195, 59.195, 59.2025, 59.2286, 59.1711, 59.1777, 59.1782, 59.2726, 
    59.2347, 59.2055, 59.2022, 59.1695, 59.1671, 59.1706, 59.1745, 59.1649, 
    59.177, 59.1717, 59.1746, 59.1647, 59.1843, 59.1803, 59.1835, 59.135, 
    59.128, 59.1281, 59.1339, 59.1285, 59.1344, 59.1341, 59.1335, 59.1322, 
    59.1263, 59.137, 59.1371, 59.1281, 59.1424, 59.1373, 59.1363, 59.1371, 
    59.1383, 59.16, 59.1589, 59.1585, 59.1717, 59.1858, 59.1522, 59.1539, 
    59.1686, 59.1797, 59.1815, 59.1861, 59.1828, 59.1349, 59.137, 59.1357, 
    59.1259, 59.1313, 59.1338, 59.1352, 59.1347, 59.135, 59.1371, 59.1353, 
    59.1354, 59.1338, 59.1706, 59.1752, 59.1742, 59.1764, 59.1767, 59.1944, 
    59.1885, 59.1733, 59.1801, 59.1754, 59.1844, 59.1929, 59.1805, 59.1937, 
    59.1704, 59.177, 59.1735, 59.1736, 59.1751, 59.1794, 59.1794, 59.1752, 
    59.1754, 59.1815, 59.1768, 59.1936, 59.192, 59.1934, 59.1934, 59.194, 
    59.1907, 59.1943, 59.1934, 59.1923, 59.1931, 59.1922, 59.1929, 59.1934, 
    59.1932, 59.1933, 59.1933, 59.1932, 59.1932, 59.1863, 59.1932, 59.1892, 
    59.1934, 59.1936, 59.194, 59.1914, 59.1909, 59.1909, 59.193, 59.1937, 
    59.1943, 50.6209, 66.8307, 59.1983, 59.1961, 59.1965, 58.6559, 58.6522, 
    58.6348, 59.2002, 58.9037, 50.8049, 59.1976, 59.1986, 59.1801, 59.202, 
    59.247, 59.201, 59.2048, 59.2051, 59.2041, 59.1933, 59.1933, 59.2007, 
    59.2041, 59.2076, 59.2099, 59.1639, 59.1604, 59.1615, 59.1208, 59.1162, 
    59.0958, 59.0947, 59.0912, 59.0917, 59.095, 59.0952, 59.0918, 59.0989, 
    59.0965, 59.0937, 59.0956, 59.0957, 59.095, 59.0949, 59.0953, 59.0961, 
    59.0936, 59.0949, 59.0972, 59.0966, 59.0998, 59.0907, 59.0932, 59.0977, 
    59.104, 59.1062, 59.1115, 59.1152, 59.1152, 59.1192, 59.1271, 59.1355, 
    59.1361, 59.1376, 59.1602, 59.1497, 59.1757, 59.1804, 59.1772, 59.1685, 
    59.1996, 59.1768, 59.188, 59.2066, 59.2089, 59.2195, 59.2212, 59.2203, 
    59.2213, 59.2237, 59.2271, 59.2255, 59.223, 59.2241, 59.2193, 59.2303, 
    59.2213, 59.2229, 59.2201, 59.2207, 59.2236, 59.2274, 59.21, 59.2098, 
    59.2113, 59.2128, 59.2162, 59.2088, 59.2075, 59.2044, 59.2086, 59.2044, 
    59.2104, 59.2086, 59.2087, 59.2087, 59.2093, 59.2077, 59.2096, 59.2096, 
    59.1941, 59.1853, 59.1878, 59.1883, 59.1789, 59.1864, 59.1845, 59.1818, 
    59.1648, 59.1617, 59.1749, 59.1647, 59.1664, 59.1847, 59.1872, 59.1316, 
    59.1415, 59.1414, 59.1509, 59.1833, 59.1959, 59.1956, 59.1957, 59.1986, 
    59.1978, 59.1987, 59.2005, 59.201, 59.1981, 59.2005, 59.1928, 59.193, 
    59.1905, 59.2066, 59.2032, 59.204, 59.1981, 59.2025, 59.1991, 59.1985, 
    59.198, 59.1978, 59.1928, 59.1958, 59.1945, 59.1968, 59.2036, 59.1974, 
    59.1984, 59.1982, 59.185, 59.1874, 59.1773, 59.1856, 59.1845, 59.1904, 
    59.1875, 59.1856, 59.1821, 59.1795, 59.166, 59.1428, 59.1279, 59.12, 
    59.1236, 59.1215, 59.1008, 59.0901, 59.0876, 59.0749, 59.0959, 59.093, 
    59.0899, 59.0953, 59.0939, 59.0939, 59.1069, 59.1092, 59.1169, 59.1183, 
    59.1254, 59.1114, 59.164, 59.1638, 59.1565, 59.1684, 59.1759, 59.1755, 
    59.1567, 59.1356, 59.1636, 59.1356, 59.1607, 59.134, 59.1343, 59.1344, 
    59.1725, 59.1724, 59.2042, 59.2165, 59.2139, 59.209, 59.2094, 59.208, 
    59.2224, 59.2049, 59.22, 59.2135, 59.2072, 59.2111, 59.2861, 59.2137, 
    59.2, 59.2029, 59.2065, 59.2081, 59.2032, 59.2073, 59.2144, 59.2194, 
    59.2026, 59.2067, 59.2178, 59.2138, 59.2142, 59.2117, 59.2082, 59.2053, 
    59.214, 59.2135, 59.2142, 59.2119, 59.2122, 59.212, 59.205, 59.1959, 
    59.219, 59.214, 59.2184, 59.2099, 59.2123, 59.1802, 59.1884, 59.2107, 
    59.015, 59.0241, 59.2285, 59.2268, 59.2359, 59.2096, 59.2085, 59.2, 
    59.1999, 59.2033, 59.2071, 59.2096, 59.1891, 59.1887, 59.177, 59.1889, 
    59.2, 59.2075, 59.1893, 59.1889, 59.1788, 59.1811, 59.1805, 59.1852, 
    59.1379, 59.1393, 59.1431, 59.1349, 59.1349, 59.133, 59.1364, 59.1366, 
    59.1118, 59.1256, 59.1955, 59.1998, 59.1356, 59.1511, 59.1868, 59.1994, 
    59.2002, 59.2003, 59.1936, 59.1976, 59.1974, 59.1936, 59.194, 59.1943, 
    59.2124, 59.2155, 59.1825, 59.19, 59.1831, 59.1884, 59.1806, 59.1882, 
    59.1745, 59.1524, 59.1659, 59.1522, 59.1621, 59.1839, 59.1794, 59.2095, 
    59.054, 59.1836, 59.174, 59.1737, 59.1974, 59.1821, 59.1701, 59.1786, 
    59.1791, 59.1951, 59.197, 59.1891, 59.1865, 59.1917, 59.1905, 59.1892, 
    59.2082, 59.1832, 59.1642, 59.1806, 59.1661, 59.1828, 59.1987, 59.1982, 
    59.1947, 59.2141, 59.146, 59.1314, 59.0937, 59.0854, 59.1165, 59.1177, 
    59.1182, 59.1103, 59.1104, 59.1411, 59.1572, 59.162, 59.1691, 59.1758, 
    59.181, 59.1789, 59.1842, 59.1891, 59.1883, 59.1851, 59.1875, 59.2029, 
    59.1868, 59.1893, 59.1972, 59.1979, 59.1972, 59.2566, 59.1898, 59.172, 
    59.1458, 59.146, 59.1332, 59.1342, 59.1366, 59.1367, 59.1331, 59.1346, 
    59.1281, 59.1098, 59.1099, 59.1336, 59.1339, 59.1273, 59.1189, 59.1166, 
    59.1176, 59.12, 59.1373, 59.1382, 59.1398, 59.1533, 59.1573, 59.1618, 
    59.1605, 59.1625, 59.194, 59.2001, 59.1874, 59.1777, 59.1768, 59.1772, 
    59.1664, 59.1632, 59.162, 59.17, 59.1827, 59.1748, 59.1857, 59.1913, 
    59.1767, 59.1964, 59.2054, 59.2067, 59.2052, 59.2021, 59.2001, 59.2015, 
    59.2021, 59.1967, 59.1964, 59.1964, 59.1964, 59.1969, 59.1967, 59.2021, 
    59.2007, 59.2014, 59.1937, 59.2015, 59.193, 59.1923, 59.1903, 59.1912, 
    59.2048, 59.2048, 59.1872, 59.1777, 59.1868, 59.1737, 59.1707, 59.1526, 
    59.1673, 59.168, 59.1726, 59.176, 59.1676, 59.1527, 59.1399, 59.1409, 
    59.124, 59.1343, 59.1309, 59.1317, 59.1326, 59.1371, 59.1184, 59.0616, 
    59.1219, 59.137, 59.1371, 59.1256, 59.138, 59.1445, 59.1372, 59.1339, 
    59.1503, 59.1495, 59.1354, 59.1311, 59.1356, 59.1337, 59.1434, 59.1482, 
    59.141, 59.1489, 59.1465, 59.1447, 59.1523, 59.1551, 59.1552, 59.1401, 
    59.139, 59.1472, 59.1463, 59.174, 59.1613, 59.1782, 59.1772, 59.1102, 
    59.0936, 59.0941, 59.0947, 59.0955, 59.0955, 59.0723, 59.0957, 59.1168, 
    59.1173, 59.1209, 59.1299, 59.1287, 59.1519, 59.1516, 59.1611, 59.1611, 
    59.1846, 59.1654, 59.1726, 59.1805, 59.2381, 59.2353, 59.1862, 59.1827, 
    59.2823, 59.1778, 59.1785, 59.1777, 59.204, 59.2018, 59.2036, 59.1989, 
    59.199, 59.1975, 59.1978, 59.1965, 59.1983, 59.1981, 59.1968, 59.199, 
    59.2077, 59.205, 59.2025, 59.2066, 59.2029, 59.202, 59.1987, 59.1995, 
    59.1982, 59.1944, 59.2006, 59.2223, 59.1911, 59.1897, 59.191, 59.1895, 
    59.1838, 59.1815, 59.1896, 59.1894, 59.1759, 59.1772, 59.1906, 59.2144, 
    59.1908, 59.1764, 59.1347, 59.1607, 59.1387, 59.1449, 59.1428, 59.1374, 
    59.136, 59.134, 59.1922, 59.1706, 59.137, 59.1363, 59.1256, 59.1171, 
    59.1064, 59.1122, 59.1321, 59.1357, 59.1258, 59.1367, 59.1239, 59.1255, 
    59.1278, 59.1362, 59.1286, 59.1321, 59.1579, 59.1321, 59.099, 59.1107, 
    59.0947, 59.0951, 59.0952, 59.0962, 59.0927, 59.0962, 59.0937, 59.0929, 
    59.0463, 59.0506, 59.1078, 59.1174, 59.1173, 59.1642, 59.0955, 59.1335, 
    59.1359, 59.1397, 59.1359, 59.1374, 59.1359, 59.1339, 59.1359, 59.1347, 
    59.1358, 59.134, 59.134, 59.1244, 59.1352, 59.1343, 59.1356, 59.1338, 
    59.1401, 59.1416, 59.1363, 59.1356, 59.1359, 59.1448, 59.1346, 59.136, 
    59.135, 59.1318, 59.1331, 59.1334, 59.1363, 59.1367, 59.118, 59.1343, 
    59.1339, 59.142, 59.1427, 59.1419, 59.1316, 59.1411, 59.1168, 59.1238, 
    59.1278, 59.1146, 59.1088, 59.1054, 59.0976, 59.1464, 59.1947, 59.2026, 
    59.2031, 59.2027, 59.2144, 59.1852, 59.1898, 59.1903, 59.1889, 59.1859, 
    59.1822, 59.1892, 59.1992, 59.178, 59.1673, 59.1927, 59.1775, 59.1856, 
    59.1856, 59.1973, 59.1828, 59.1716, 59.1818, 59.1692, 59.1921, 59.1864, 
    59.1622, 59.1587, 59.1547, 59.1539, 59.1556, 59.1629, 59.0973, 59.0945, 
    59.1097, 59.1032, 59.0949, 59.087, 59.0916, 59.0937, 59.0955, 59.0107, 
    59.0957, 59.1, 59.1017, 59.12, 59.1192, 59.1184, 59.1153, 59.1329, 
    59.1329, 59.1311, 59.1303, 59.1562, 59.1563, 59.1557, 59.1562, 59.1551, 
    59.1585, 59.1708, 59.1632, 59.162, 59.1637, 59.1676, 59.1678, 59.1589, 
    59.163, 59.1637, 59.1653, 59.1669, 59.1656, 59.1581, 59.136, 59.1456, 
    59.1481, 59.1478, 59.1371, 59.1454, 59.1242, 59.1336, 59.1356, 59.1278, 
    59.1343, 59.1372, 59.1358, 59.14, 59.1343, 59.1334, 59.1344, 59.1352, 
    59.1507, 59.1525, 59.1521, 59.1527, 59.1694, 59.1619, 59.1575, 59.1526, 
    59.1634, 59.1546, 59.1584, 59.1565, 59.1402, 59.1172, 59.0966, 59.0924, 
    59.0938, 59.0949, 59.0739, 59.1183, 59.1196, 59.1185, 59.1199, 59.1272, 
    59.1376, 59.1317, 59.1564, 59.1368, 59.1819, 59.2124, 59.1848, 59.1396, 
    59.1359, 59.1356, 59.1406, 59.1357, 59.1394, 59.1356, 59.1357, 59.1325, 
    59.1351, 59.1308, 59.1304, 59.1302, 59.1243, 59.1264, 59.1308, 59.1309, 
    59.1329, 59.1236, 59.1318, 59.1324, 59.1307, 59.1304, 59.1302, 59.1568, 
    59.1602, 59.1624, 59.1536, 59.1592, 59.1699, 59.1685, 59.1893, 59.0942, 
    59.0951, 59.0976, 59.0892, 59.0858, 59.0935, 59.0879, 59.0942, 59.0919, 
    59.0935, 59.0948, 59.1026, 59.096, 59.0955, 59.0956, 59.096, 59.0948, 
    59.0898, 59.0926, 59.0933, 59.1044, 59.1261, 59.1231, 59.123, 59.1195, 
    59.1241 ;

 location_class = "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", 
    "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", 
    "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", 
    "G", "G", "G", "G", "2", "2", "A", "A", "2", "1", "3", "3", "B", "G", 
    "G", "G", "G", "G", "G", "G", "B", "G", "G", "B", "G", "B", "G", "G", 
    "B", "B", "B", "B", "G", "B", "B", "G", "B", "G", "B", "A", "B", "G", 
    "G", "B", "G", "G", "B", "G", "G", "B", "G", "B", "1", "B", "B", "B", 
    "B", "B", "B", "B", "G", "G", "G", "0", "G", "B", "G", "B", "B", "B", 
    "B", "B", "B", "2", "1", "1", "B", "B", "B", "B", "B", "B", "B", "B", 
    "B", "B", "B", "A", "3", "B", "B", "1", "B", "B", "B", "B", "B", "B", 
    "G", "B", "B", "B", "2", "B", "B", "1", "0", "A", "1", "G", "2", "2", 
    "3", "2", "1", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", 
    "2", "2", "A", "B", "G", "B", "2", "2", "2", "B", "B", "G", "B", "B", 
    "B", "2", "B", "3", "3", "2", "A", "2", "2", "2", "3", "2", "B", "G", 
    "G", "G", "G", "G", "G", "G", "G", "G", "G", "A", "G", "G", "G", "B", 
    "B", "B", "B", "B", "B", "B", "B", "B", "1", "B", "2", "1", "B", "B", 
    "A", "B", "G", "G", "B", "G", "G", "G", "B", "B", "A", "B", "A", "B", 
    "2", "A", "A", "2", "2", "B", "3", "2", "2", "2", "G", "A", "2", "B", 
    "0", "B", "0", "A", "B", "G", "G", "G", "G", "G", "G", "G", "G", "G", 
    "G", "B", "A", "B", "G", "G", "1", "G", "B", "B", "1", "A", "G", "1", 
    "2", "G", "1", "G", "0", "G", "3", "2", "B", "3", "B", "1", "3", "3", 
    "A", "A", "2", "G", "G", "B", "G", "G", "G", "G", "G", "G", "G", "G", 
    "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "B", 
    "G", "0", "B", "B", "B", "2", "G", "B", "A", "B", "1", "A", "3", "B", 
    "A", "1", "B", "B", "A", "B", "G", "B", "B", "G", "G", "G", "G", "G", 
    "G", "G", "G", "G", "G", "2", "3", "2", "B", "3", "3", "B", "1", "A", 
    "B", "3", "3", "3", "B", "3", "2", "A", "2", "B", "3", "3", "B", "2", 
    "1", "B", "B", "A", "A", "B", "B", "B", "B", "B", "B", "3", "B", "G", 
    "0", "G", "G", "A", "B", "2", "G", "2", "G", "1", "A", "A", "B", "2", 
    "A", "G", "1", "G", "1", "G", "A", "G", "A", "B", "G", "G", "G", "G", 
    "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "B", "B", 
    "G", "G", "G", "B", "B", "G", "G", "G", "G", "B", "G", "B", "A", "G", 
    "A", "B", "G", "A", "3", "G", "B", "B", "B", "B", "B", "B", "G", "0", 
    "B", "B", "G", "B", "B", "B", "G", "G", "G", "G", "G", "G", "G", "B", 
    "G", "B", "G", "B", "B", "A", "A", "B", "B", "B", "B", "B", "A", "G", 
    "G", "G", "G", "B", "G", "G", "2", "G", "0", "G", "B", "G", "B", "1", 
    "1", "B", "B", "B", "G", "1", "1", "1", "2", "A", "1", "2", "2", "3", 
    "B", "G", "G", "B", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", 
    "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", 
    "2", "B", "G", "B", "G", "B", "G", "B", "A", "G", "B", "B", "A", "B", 
    "B", "B", "3", "G", "G", "G", "1", "B", "G", "G", "1", "G", "2", "G", 
    "2", "B", "A", "0", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", 
    "G", "G", "B", "B", "B", "B", "G", "B", "B", "G", "B", "B", "A", "A", 
    "A", "B", "B", "B", "3", "G", "G", "B", "B", "A", "B", "3", "3", "B", 
    "B", "B", "G", "3", "1", "B", "1", "B", "B", "B", "B", "B", "B", "1", 
    "B", "1", "B", "B", "B", "B", "G", "G", "G", "B", "B", "G", "0", "B", 
    "B", "B", "1", "1", "1", "G", "3", "3", "A", "B", "3", "B", "1", "B", 
    "1", "2", "1", "G", "B", "B", "B", "G", "G", "G", "G", "G", "G", "G", 
    "G", "A", "G", "G", "G", "G", "G", "B", "G", "G", "G", "B", "G", "B", 
    "B", "G", "G", "G", "B", "B", "B", "2", "G", "B", "B", "G", "B", "0", 
    "G", "B", "G", "B", "2", "G", "G", "G", "G", "1", "0", "G", "B", "G", 
    "1", "G", "G", "G", "G", "2", "G", "B", "G", "G", "G", "G", "A", "1", 
    "2", "B", "1", "3", "3", "3", "2", "3", "3", "A", "1", "1", "2", "2", 
    "A", "1", "3", "2", "3", "B", "B", "A", "G", "G", "G", "G", "G", "G", 
    "G", "G", "G", "G", "B", "B", "B", "G", "G", "B", "G", "0", "2", "3", 
    "0", "2", "3", "A", "2", "3", "3", "B", "3", "B", "2", "3", "B", "B", 
    "B", "G", "G", "G", "G", "G", "G", "G", "B", "B", "B", "B", "1", "B", 
    "A", "B", "A", "A", "B", "A", "2", "1", "A", "G", "A", "B", "G", "G", 
    "G", "G", "B", "B", "G", "B", "G", "B", "B", "2", "0", "1", "A", "2", 
    "B", "A", "3", "3", "B", "A", "3", "B", "B", "B", "G", "G", "1", "G", 
    "G", "B", "B", "B", "B", "2", "A", "A", "B", "B", "B", "B", "1", "1", 
    "B", "2", "B", "A", "A", "G", "G", "G", "G", "0", "B", "B", "B", "B", 
    "B", "B", "G", "G", "B", "B", "B", "G", "B", "G", "G", "B", "B", "B", 
    "B", "G", "B", "B", "G", "B", "B", "G", "3", "1", "A", "3", "B", "B", 
    "A", "B", "G", "G", "B", "3", "2", "B", "A", "A", "G", "2", "A", "B", 
    "A", "2", "B", "B", "B", "B", "B", "B", "B", "B", "B", "G", "G", "B", 
    "G", "G", "G", "G", "G", "G", "0", "B", "G", "1", "2", "B", "G", "A", 
    "1", "B", "1", "1", "3", "2", "G", "A", "1", "2", "2", "3", "1", "3", 
    "A", "A", "1", "B", "B", "G", "G", "G", "G", "G", "G", "G", "G", "G", 
    "G", "G", "G", "G", "G", "2", "1", "B", "2", "B", "B", "3", "B", "2", 
    "3", "B", "3", "B", "B", "2", "3", "2", "1", "B", "B", "1", "A", "0", 
    "B", "B", "B", "B", "G", "G", "G", "G", "G", "G", "G", "G", "2", "B", 
    "G", "G", "G", "G", "A", "A", "B", "B", "B", "B", "B", "B", "B", "B", 
    "B", "A", "B", "G", "B", "G", "B", "G", "G", "B", "A", "B", "B", "G", 
    "B", "G", "A", "B", "B", "A", "B", "A", "A", "B", "A", "1", "B", "1", 
    "1", "3", "B", "B", "G", "B", "1", "G", "G", "1", "B", "B", "1", "B", 
    "B", "B", "1", "2", "A", "B", "A", "A", "A", "B", "2", "2", "2", "G", 
    "1", "G", "0", "G", "2", "G", "3", "G", "2", "B", "G", "G", "G", "G", 
    "G", "B", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", 
    "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "A", 
    "G", "B", "G", "G", "A", "B", "B", "G", "G", "2", "1", "3", "2", "G", 
    "2", "3", "G", "G", "2", "3", "G", "G", "2", "G", "1", "G", "2", "3", 
    "G", "A", "G", "A", "G", "3", "G", "A", "G", "B", "B", "B", "B", "B", 
    "G", "G", "G", "G", "G", "G", "G", "B", "B", "B", "B", "B", "A", "0", 
    "3", "1", "3", "2", "1", "G", "B", "2", "B", "0", "2", "3", "B", "B", 
    "G", "B", "G", "B", "B", "B", "B", "B", "G", "G", "B", "G", "G", "B", 
    "B", "A", "B", "B", "G", "B", "1", "G", "B", "B", "G", "B", "G", "B", 
    "G", "G", "G", "G", "B", "G", "G", "G", "G", "2", "0", "1", "1", "B", 
    "3", "B", "3", "B", "3", "3", "2", "B", "1", "3", "G", "B", "G", "G", 
    "A", "G", "B", "G", "G", "G", "G", "G", "B", "A", "B", "G", "G", "G", 
    "G", "G", "G", "B", "B", "A", "G", "A", "G", "B", "G", "G", "G", "3", 
    "3", "3", "A", "3", "2", "2", "3", "3", "3", "G", "1", "3", "0", "3", 
    "3", "B", "G", "G", "B", "G", "G", "G", "B", "G", "G", "1", "2", "2", 
    "A", "B", "1", "3", "2", "B", "2", "3", "3", "B", "1", "1", "2", "3", 
    "A", "B", "A", "B", "B", "0", "G", "B", "B", "G", "B", "B", "A", "3", 
    "B", "G", "B", "G", "G", "B", "B", "B", "B", "G", "G", "G", "G", "G", 
    "B", "1", "G", "G", "G", "G", "B", "G", "G", "B", "G", "G", "G", "3", 
    "B", "G", "A", "G", "B", "B", "A", "1", "B", "B", "B", "G", "B", "2", 
    "G", "G", "B", "G", "B", "G", "B", "G", "G", "G", "G", "G", "B", "G", 
    "A", "G", "G", "2", "B", "G", "G", "2", "2", "2", "1", "3", "1", "2", 
    "1", "1", "A", "1", "1", "1", "1", "1", "1", "A", "B", "A", "1", "A", 
    "G", "2", "1", "A", "B", "2", "B", "A", "2", "0", "B", "B", "B", "G", 
    "B", "A", "A", "B", "B", "B", "B", "2", "0", "B", "G", "B", "B", "B", 
    "G", "G", "G", "B", "B", "G", "3", "1", "1", "2", "1", "B", "B", "2", 
    "0", "G", "G", "B", "B", "G", "2", "B", "B", "G", "G", "B", "B", "1", 
    "G", "B", "B", "B", "G", "B", "G", "B", "B", "B", "A", "B", "B", "A", 
    "B", "B", "1", "1", "B", "G", "B", "B", "B", "1", "B", "B", "0", "A", 
    "A", "A", "B", "A", "B", "3", "2", "A", "1", "B", "G", "G", "G", "G", 
    "G", "G", "B", "G", "G", "G", "G", "B", "B", "A", "B", "B", "B", "B", 
    "G", "G", "A", "B", "B", "2", "A", "A", "3", "B", "B", "B", "G", "G", 
    "G", "1", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", 
    "1", "B", "G", "B", "3", "1", "A", "A", "B", "B", "B", "A", "B", "A", 
    "B", "3", "3", "3", "B", "3", "B", "G", "G", "B", "B", "B", "B", "B", 
    "B", "B", "B", "B", "B", "A", "1", "2", "2", "B", "2", "1", "B", "G", 
    "G", "G", "G", "G", "G", "B", "G", "2", "B", "B", "G", "G", "G", "G", 
    "G", "G", "G", "G", "G", "G", "G", "G", "G", "B", "3", "B", "B", "G", 
    "3", "1", "B", "B", "B", "B", "1", "G", "1", "B", "G", "B", "G", "B", 
    "B", "G", "B", "B", "G", "G", "A", "B", "G", "A", "B", "B", "G", "G", 
    "G", "B", "B", "B", "B", "B", "G", "B", "B", "G", "B", "B", "B", "G", 
    "G", "G", "3", "B", "B", "1", "B", "B", "B", "3", "2", "B", "2", "3", 
    "2", "3", "3", "3", "A", "1", "A", "2", "1", "3", "B", "G", "B", "G", 
    "G", "G", "G", "1", "G", "G", "B", "G", "A", "B", "B", "B", "B", "B", 
    "B", "A", "G", "B", "B", "B", "B", "B", "B", "G", "G", "2", "1", "G", 
    "B", "G", "G", "B", "B", "B", "A", "B", "B", "G", "G", "G", "G", "G", 
    "B", "2", "B", "B", "3", "B", "A", "2", "A", "2", "2", "B", "B", "3", 
    "A", "B", "0", "G", "B", "2", "B", "B", "B", "B", "A", "G", "G", "G", 
    "G", "G", "G", "G", "G", "G", "G", "B", "B", "A", "G", "B", "G", "B", 
    "B", "A", "B", "1", "A", "A", "G", "1", "0", "B", "0", "B", "A", "1", 
    "2", "G", "2", "1", "1", "3", "B", "B", "G", "G", "G", "0", "G", "B", 
    "B", "B", "B", "B", "B", "B", "B", "G", "B", "G", "G", "G", "G", "B", 
    "B", "B", "G", "G", "G", "G", "G", "A", "B", "G", "B", "G", "A", "B", 
    "B", "G", "B", "B", "B", "A", "B", "B", "1", "A", "G", "B", "1", "2", 
    "1", "B", "B", "B", "B", "G", "3", "A", "1", "G", "B", "B", "3", "A", 
    "B", "A", "B", "1", "B", "2", "A", "B", "B", "B", "B", "B", "3", "B", 
    "1", "G", "G", "B", "3", "B", "A", "G", "B", "A", "B", "B", "A", "3", 
    "A", "3", "1", "3", "2", "B", "0", "2", "3", "0", "A", "B", "1", "G", 
    "G", "G", "B", "G", "B", "B", "A", "B", "G", "B", "B", "B", "B", "G", 
    "G", "B", "B", "G", "A", "A", "B", "B", "B", "1", "G", "B", "G", "B", 
    "G", "A", "G", "B", "A", "2", "B", "2", "G", "G", "G", "G", "G", "G", 
    "B", "G", "B", "G", "B", "B", "G", "G", "B", "G", "A", "A", "2", "3", 
    "G", "A", "B", "B", "A", "B", "3", "G", "1", "G", "G", "A", "B", "B", 
    "B", "A", "A", "B", "B", "B", "2", "B", "3", "B", "G", "G", "G", "G", 
    "G", "G", "G", "G", "G", "G", "G", "B", "B", "G", "A", "B", "G", "A", 
    "B", "3", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "A", "G", 
    "G", "B", "G", "B", "B", "G", "B", "G", "B", "G", "B", "B", "B", "G", 
    "1", "G", "A", "G", "B", "G", "G", "A", "A", "B", "3", "A", "B", "B", 
    "B", "G", "B", "G", "G", "A", "1", "2", "B", "A", "G", "B", "G", "A", 
    "2", "B", "A", "B", "3", "B", "B", "A", "A", "A", "A", "B", "B", "B", 
    "B", "G", "G", "B", "3", "B", "B", "1", "B", "B", "B", "G", "B", "B", 
    "G", "A", "A", "B", "A", "B", "B", "1", "2", "A", "G", "0", "A", "G", 
    "B", "B", "B", "G", "B", "2", "G", "G", "G", "G", "A", "G", "A", "G", 
    "B", "G", "B", "B", "A", "B", "B", "G", "0", "1", "1", "B", "B", "A", 
    "0", "A", "A", "2", "B", "B", "B", "B", "B", "G", "G", "G", "G", "G", 
    "A", "G", "B", "1", "B", "B", "G", "G", "G", "G", "G", "G", "G", "B", 
    "B", "B", "2", "A", "1", "B", "A", "G", "B", "3", "3", "A", "3", "B", 
    "A", "2", "B", "A", "G", "G", "B", "B", "B", "G", "G", "G", "G", "G", 
    "A", "B", "B", "A", "G", "B", "B", "3", "1", "B", "1", "B", "2", "2", 
    "2", "2", "2", "G", "G", "B", "1", "3", "0", "A", "B", "A", "A", "2", 
    "G", "G", "G", "G", "G", "G", "0", "B", "A", "2", "B", "0", "B", "1", 
    "B", "A", "B", "A", "B", "B", "G", "B", "G", "B", "G", "A", "G", "G", 
    "G", "G", "G", "G", "G", "G", "B", "B", "B", "B", "G", "G", "G", "B", 
    "0", "A", "B", "B", "B", "G", "G", "G", "G", "0", "2", "B", "G", "B", 
    "B", "B", "G", "G", "3", "1", "B", "B", "G", "A", "A", "A", "G", "A", 
    "B", "G", "G", "B", "1", "B", "B", "A", "G", "G", "G", "G", "A", "B", 
    "G", "A", "B", "B", "B", "B", "G", "B", "B", "B", "B", "B", "B", "A", 
    "1", "2", "1", "2", "3", "3", "3", "G", "A", "A", "G", "G", "G", "B", 
    "G", "G", "G", "B", "G", "B", "G", "A", "G", "G", "G", "G", "B", "B", 
    "G", "B", "G", "0", "G", "G", "A", "G", "A", "B", "G", "B", "B", "G", 
    "B", "B", "B", "B", "G", "G", "B", "G", "B", "B", "B", "B", "2", "B", 
    "B", "1", "1", "B", "B", "0", "G", "A", "G", "B", "0", "2", "G", "G", 
    "B", "B", "G", "B", "B", "G", "G", "G", "B", "B", "B", "A", "B", "G", 
    "G", "G", "G", "G", "G", "B", "B", "A", "1", "1", "B", "A", "2", "2", 
    "A", "B", "B", "2", "0", "1", "0", "1", "G", "A", "A", "2", "2", "3", 
    "3", "B", "A", "G", "G", "G", "B", "3", "B", "3", "2", "B", "B", "G", 
    "G", "3", "3", "A", "2", "3", "B", "3", "A", "1", "3", "B", "B", "A", 
    "G", "G", "A", "2", "G", "B", "A", "G", "A", "B", "G", "B", "B", "B", 
    "B", "A", "B", "B", "B", "G", "B", "G", "G", "G", "B", "B", "0", "B", 
    "B", "B", "G", "B", "B", "A", "B", "A", "B", "3", "G", "2", "A", "2", 
    "G", "B", "1", "B", "3", "G", "3", "1", "A", "G", "A", "1", "B", "B", 
    "G", "G", "G", "G", "B", "B", "G", "G", "G", "B", "G", "G", "B", "B", 
    "B", "1", "G", "G", "G", "B", "G", "G", "B", "G", "B", "B", "G", "B", 
    "G", "G", "B", "G", "G", "B", "A", "G", "1", "B", "G", "B", "B", "G", 
    "B", "B", "B", "B", "0", "G", "B", "G", "1", "B", "G", "A", "B", "B", 
    "B", "2", "2", "1", "2", "0", "2", "B", "G", "B", "B", "G", "B", "B", 
    "B", "G", "B", "G", "1", "G", "G", "G", "G", "G", "G", "G", "B", "2", 
    "B", "G", "G", "G", "G", "3", "1", "B", "B", "0", "G", "1", "G", "0", 
    "2", "2", "B", "2", "1", "1", "1", "1", "B", "B", "3", "2", "3", "1", 
    "1", "B", "G", "G", "G", "G", "G", "G", "G", "1", "1", "1", "3", "1", 
    "1", "3", "G", "2", "2", "G", "G", "1", "A", "3", "G", "B", "0", "B", 
    "2", "B", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", 
    "B", "G", "G", "0", "B", "B", "B", "B", "B", "B", "B", "B", "A", "B", 
    "B", "B", "0", "B", "B", "A", "A", "A", "2", "B", "B", "2", "2", "3", 
    "B", "A", "B", "2", "3", "2", "3", "2", "2", "B", "2", "B", "A", "2", 
    "1", "2", "3", "A", "0", "1", "2", "B", "B", "G", "G", "G", "G", "G", 
    "G", "G", "G", "G", "G", "1", "2", "A", "3", "2", "B", "1", "G", "B", 
    "A", "1", "B", "B", "B", "A", "B", "B", "B", "A", "A", "G", "3", "G", 
    "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "B", "B", 
    "G", "G", "B", "G", "G", "B", "B", "B", "A", "B", "B", "A", "B", "1", 
    "3", "B", "3", "B", "1", "A", "2", "1", "B", "3", "B", "1", "2", "G", 
    "B", "B", "G", "G", "G", "G", "G", "G", "B", "G", "B", "G", "B", "B", 
    "A", "B", "G", "B", "0", "G", "B", "B", "G", "B", "G", "B", "G", "B", 
    "G", "B", "0", "0", "G", "B", "B", "B", "B", "B", "B", "G", "G", "G", 
    "G", "G", "B", "G", "G", "B", "B", "G", "G", "B", "1", "A", "A", "B", 
    "1", "B", "3", "B", "B", "B", "B", "B", "G", "G", "G", "G", "G", "G", 
    "G", "B", "B", "G", "G", "2", "2", "3", "A", "B", "A", "G", "B", "B", 
    "B", "B", "B", "G", "B", "G", "B", "G", "G", "A", "B", "G", "B", "B", 
    "G", "G", "G", "G", "B", "3", "2", "1", "2", "B", "3", "2", "3", "3", 
    "A", "3", "3", "3", "3", "3", "B", "A", "3", "3", "B", "B", "B", "2", 
    "B", "G", "G", "G", "2", "G", "2", "G", "B", "B", "B", "1", "A", "0", 
    "A", "G", "B", "A", "A", "B", "B", "B", "G", "0", "B", "1", "1", "B", 
    "B", "B", "A", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "B", 
    "B", "G", "2", "1", "0", "2", "G", "1", "1", "G", "B", "B", "B", "B", 
    "1", "A", "B", "1", "G", "B", "1", "G", "A", "B", "G", "G", "G", "G", 
    "G", "G", "G", "G", "G", "B", "2", "B", "1", "G", "2", "G", "B", "G", 
    "B", "B", "B", "G", "B", "B", "B", "G", "A", "A", "B", "B", "B", "A", 
    "A", "1", "G", "B", "G", "2", "B", "B", "B", "B", "G", "B", "G", "G", 
    "G", "G", "G", "B", "G", "B", "G", "G", "G", "G", "G", "G", "G", "G", 
    "G", "B", "2", "3", "B", "B", "3", "G", "3", "G", "G", "A", "B", "B", 
    "A", "G", "G", "B", "3", "G", "2", "0", "G", "G", "A", "G", "B", "B", 
    "B", "B", "1", "B", "B", "G", "G", "B", "B", "A", "B", "B", "B", "0", 
    "A", "1", "G", "B", "G", "G", "B", "B", "A", "A", "3", "B", "A", "2", 
    "B", "2", "3", "B", "A", "B", "B", "G", "B", "G", "B", "B", "G", "G", 
    "G", "B", "B", "B", "1", "A", "B", "1", "A", "B", "2", "B", "B", "B", 
    "B", "B", "B", "B", "B", "B", "G", "B", "B", "A", "B", "B", "G", "G", 
    "G", "G", "G", "G", "G", "G", "B", "B", "G", "B", "G", "G", "G", "B", 
    "B", "B", "B", "G", "B", "B", "B", "A", "B", "B", "A", "B", "2", "B", 
    "B", "B", "B", "G", "G", "B", "A", "B", "3", "G", "B", "B", "G", "G", 
    "B", "A", "A", "B", "B", "B", "B", "2", "B", "2", "G", "2", "1", "3", 
    "B", "A", "2", "1", "3", "B", "1", "B", "1", "B", "B", "2", "A", "3", 
    "G", "G", "G", "G", "G", "G", "B", "B", "B", "G", "G", "A", "0", "G", 
    "G", "B", "B", "B", "A", "G", "1", "G", "G", "B", "G", "0", "1", "G", 
    "2", "B", "G", "1", "G", "2", "B", "G", "G", "G", "G", "G", "G", "G", 
    "G", "G", "B", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", 
    "G", "G", "G", "G", "B", "B", "G", "G", "1", "G", "B", "G", "3", "2", 
    "B", "B", "B", "B", "B", "B", "A", "A", "B", "B", "B", "G", "B", "A", 
    "3", "B", "A", "G", "1", "G", "G", "3", "G", "3", "1", "2", "1", "1", 
    "1", "1", "2", "B", "A", "G", "B", "3", "B", "B", "G", "G", "B", "B", 
    "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", 
    "G", "1", "G", "G", "1", "B", "A", "B", "B", "B", "B", "B", "B", "B", 
    "B", "2", "1", "2", "1", "B", "B", "1", "G", "A", "G", "G", "G", "G", 
    "2", "0", "2", "B", "A", "B", "3", "1", "G", "1", "1", "3", "3", "G", 
    "G", "3", "3", "1", "G", "3", "G", "G", "B", "A", "B", "B", "A", "B", 
    "1", "G", "1", "G", "G", "1", "2", "G", "G", "1", "G", "B", "2", "A", 
    "B", "3", "3", "3", "3", "A", "B", "3", "A", "3", "B", "B", "1", "G", 
    "1", "B", "B", "G", "B", "B", "2", "3", "2", "A", "B", "B", "B", "B", 
    "G", "G", "B", "G", "B", "B", "G", "B", "A", "A", "G", "B", "G", "B", 
    "B", "B", "A", "B", "B", "B", "B", "A", "A", "2", "2", "B", "B", "B", 
    "B", "A", "B", "B", "B", "B", "A", "3", "3", "B", "2", "B", "G", "G", 
    "A", "B", "A", "A", "A", "B", "G", "G", "G", "B", "A", "B", "2", "2", 
    "1", "A", "B", "B", "B", "B", "2", "3", "B", "B", "B", "3", "G", "B", 
    "A", "A", "A", "3", "B", "B", "2", "B", "B", "B", "G", "1", "G", "G", 
    "G", "B", "B", "B", "B", "G", "A", "G", "1", "G", "A", "B", "A", "G", 
    "B", "1", "B", "B", "B", "B", "B", "B", "B", "G", "G", "G", "B", "G", 
    "G", "B", "G", "G", "G", "G", "B", "1", "B", "B", "G", "3", "B", "A", 
    "B", "B", "G", "G", "B", "0", "B", "1", "B", "2", "B", "B", "G", "B", 
    "B", "2", "A", "A", "0", "B", "B", "3", "A", "B", "B", "B", "B", "B", 
    "B", "B", "B", "B", "B", "G", "G", "G", "G", "B", "A", "1", "1", "3", 
    "3", "G", "G", "G", "G", "B", "B", "B", "B", "2", "1", "B", "A", "A", 
    "A", "2", "G", "0", "1", "2", "B", "1", "1", "3", "1", "A", "G", "2", 
    "2", "A", "G", "B", "G", "B", "B", "G", "G", "G", "G", "G", "G", "G", 
    "G", "G", "G", "G", "G", "G", "B", "G", "G", "G", "A", "G", "B", "G", 
    "1", "B", "G", "B", "2", "0", "3", "B", "B", "B", "3", "B", "3", "A", 
    "3", "2", "3", "1", "3", "B", "3", "A", "1", "G", "G", "G", "G", "B", 
    "G", "2", "G", "B", "B", "2", "2", "2", "3", "3", "0", "B", "3", "3", 
    "A", "A", "0", "B", "3", "A", "B", "1", "3", "B", "G", "G", "G", "G", 
    "G", "G", "G", "G", "A", "G", "B", "G", "B", "B", "G", "G", "B", "B", 
    "2", "G", "G", "A", "1", "G", "B", "G", "0", "2", "1", "G", "B", "G", 
    "A", "3", "1", "B", "B", "G", "B", "G", "B", "G", "G", "A", "B", "B", 
    "G", "G", "B", "G", "G", "1", "B", "G", "B", "G", "G", "B", "3", "G", 
    "G", "A", "3", "2", "G", "0", "G", "G", "0", "B", "B", "B", "B", "G", 
    "G", "G", "B", "B", "G", "0", "B", "G", "2", "3", "A", "A", "G", "A", 
    "G", "G", "G", "B", "B", "G", "B", "1", "0", "B", "G", "B", "B", "G", 
    "G", "G", "B", "B", "G", "G", "B", "G", "G", "A", "G", "1", "G", "2", 
    "G", "B", "B", "B", "B", "B", "B", "A", "B", "B", "B", "1", "B", "G", 
    "G", "G", "G", "B", "B", "G", "B", "B", "1", "G", "B", "G", "A", "G", 
    "B", "A", "0", "0", "A", "B", "3", "B", "B", "3", "G", "B", "B", "G", 
    "G", "G", "B", "G", "G", "B", "A", "1", "A", "B", "G", "G", "G", "G", 
    "G", "G", "A", "G", "B", "B", "B", "G", "G", "B", "B", "B", "B", "B", 
    "B", "B", "B", "B", "G", "B", "G", "B", "G", "G", "B", "G", "G", "B", 
    "B", "B", "B", "G", "B", "B", "3", "B", "2", "A", "G", "1", "3", "G", 
    "G", "G", "G", "G", "B", "G", "B", "G", "2", "3", "3", "B", "B", "B", 
    "B", "B", "B", "B", "G", "B", "B", "G", "1", "B", "B", "B", "B", "B", 
    "B", "A", "B", "B", "B", "1", "2", "A", "B", "2", "B", "B", "A", "B", 
    "A", "2", "B", "G", "B", "B", "A", "B", "B", "B", "B", "G", "G", "G", 
    "G", "B", "G", "G", "B", "B", "B", "A", "B", "B", "B", "B", "G", "G", 
    "G", "G", "B", "B", "G", "1", "1", "2", "3", "B", "1", "2", "3", "A", 
    "A", "1", "3", "3", "3", "2", "3", "3", "2", "1", "3", "2", "1", "1", 
    "2", "2", "2", "A", "B", "B", "G", "2", "B", "B", "0", "2", "G", "0", 
    "B", "B", "B", "B", "B", "B", "B", "B", "B", "B", "3", "B", "B", "B", 
    "G", "B", "B", "G", "B", "2", "G", "G", "0", "1", "B", "1", "A", "2", 
    "A", "2", "G", "2", "2", "2", "1", "B", "B", "3", "A", "B", "G", "0", 
    "G", "G", "G", "B", "G", "G", "G", "G", "G", "G", "G", "G", "G", "G", 
    "G", "G", "G", "G", "B", "B", "G", "0", "B", "1", "2", "A", "1", "A", 
    "1", "3", "B", "G", "3", "2", "G", "G", "3", "G", "A", "G", "2", "B", 
    "G", "B", "B", "B", "A", "G", "G", "B", "G", "B", "G", "G", "G", "G", 
    "B", "A", "B", "B", "B", "B", "B", "G", "B", "G", "A", "G", "B", "B", 
    "3", "2", "B", "G", "A", "B", "1", "B", "B", "B", "G", "G", "B", "A", 
    "B", "A", "3", "B", "B", "1", "2", "B", "1", "B", "A", "3", "B", "2", 
    "B", "B", "3", "3", "2", "2", "3", "3", "1", "B", "3", "3", "1", "B", 
    "B", "2", "1", "A", "A", "A", "G", "A", "A", "B", "B", "G", "B", "B", 
    "G", "G", "G", "G", "B", "G", "G", "B", "G", "G", "B", "G", "G", "B", 
    "G", "A", "G", "G", "G", "G", "G", "2", "B", "G", "2", "G", "G", "G", 
    "3", "A", "A", "A", "1", "G", "B", "A", "B", "B", "B", "1", "G", "G", 
    "B", "G", "G", "G", "G", "B", "B", "G", "B", "B", "G", "A", "A", "G", 
    "B", "B", "B", "A", "B", "B", "B", "B", "B", "B", "G", "G", "B", "B", 
    "G", "G", "B", "B", "A", "B", "B", "A", "B", "B", "B", "B", "G", "G", 
    "G", "B", "A", "B", "B", "2", "B", "B", "B", "B", "A", "B", "B", "3", 
    "B", "2", "B", "B", "B", "B", "B", "B", "B", "B", "B", "B", "G", "G", 
    "B", "B", "G", "G", "B", "B", "B", "0", "3", "G", "B", "B", "G", "B", 
    "G", "G", "G", "B", "2", "B", "B", "B", "B", "B", "B", "1", "B", "B", 
    "B", "B", "A", "B", "B", "B", "A", "B", "G", "B", "G", "B", "B", "G", 
    "G", "G", "0", "G", "1", "G", "G", "2", "B", "2", "G", "A", "G", "B", 
    "G", "G", "G", "G", "G", "G", "G", "B", "G", "A", "G", "B", "B", "2", 
    "B", "A", "2", "B", "B", "0", "A", "B", "B", "B", "2", "B", "B", "G", 
    "Z", "A", "B", "B", "G", "B", "B", "G", "A", "B", "B", "0", "G", "G", 
    "G", "G", "G", "G", "G", "G", "G", "G", "2", "A", "B", "B", "1", "B", 
    "A", "3", "3", "3", "3", "A", "B", "3", "B", "3", "3", "2", "3", "A", 
    "3", "2", "3", "1", "A", "G", "G", "B", "A", "A", "G", "B", "B", "B", 
    "G", "B", "G", "G", "G", "B", "B", "G", "G", "B", "B", "G", "3", "3", 
    "G", "B", "B", "B", "3", "B", "0", "A", "3", "B", "3", "B", "B", "B", 
    "3", "B", "1", "2", "3", "G", "3", "B", "A", "B", "1", "3", "B", "G", 
    "3", "A", "1", "A", "A", "2", "2", "B", "G", "B", "B", "B", "G", "G", 
    "B", "G", "G", "G", "G", "G", "G", "G", "G", "B", "2", "B", "B", "G", 
    "G", "1", "1", "B", "B", "B", "A", "B", "A", "B", "B", "B", "G", "B", 
    "B", "B", "G", "G", "A", "G", "G", "B", "A", "1", "B", "A", "B", "B", 
    "G", "G", "G", "G", "G", "G", "G", "G", "B", "G", "G", "G", "A", "B", 
    "1", "1", "A", "B", "2", "A", "A", "3", "3", "B", "A", "A", "B", "2", 
    "B", "B", "A", "B", "G", "1", "A", "B", "B", "G", "B", "G", "B", "A", 
    "3", "B", "B", "B", "0", "B", "B", "G", "3", "G", "B", "2", "B", "B", 
    "A", "1", "B", "2", "B", "B", "1", "A", "B", "1", "2", "1", "B", "2", 
    "2", "3", "2", "A", "B", "B", "1", "3", "B", "B", "B", "G", "B", "B", 
    "A", "G", "G", "G", "G", "G", "G", "G", "B", "B", "A", "G", "B", "B", 
    "B", "1", "B", "B", "B", "B", "B", "B", "B", "A", "1", "B", "A", "B", 
    "A", "B", "B", "B", "B", "1", "B", "B", "0", "B", "3", "B", "B", "B", 
    "G", "G", "B", "B", "B", "B", "B", "B", "B", "B", "A", "A", "2", "B", 
    "B", "B", "B", "0", "0", "B", "G", "B", "A", "2", "2", "1", "G", "G", 
    "G", "G", "B", "G", "G", "G", "A", "A", "B", "G", "1", "3", "A", "B", 
    "2", "A", "B", "G", "B", "B", "B", "G", "A", "B", "B", "B", "B", "B", 
    "B", "B", "3", "B", "A", "B", "B", "B", "B", "G", "G", "A", "A", "B", 
    "B", "B", "G", "B", "B", "A", "B", "B", "G", "G", "G", "G", "G", "B", 
    "G", "G", "3", "A", "A", "2", "2", "G", "G", "G", "0", "B", "B", "G", 
    "G", "B", "0", "B", "B", "B", "1", "B", "B", "B", "B", "B", "B", "B", 
    "A", "B", "G", "1", "G", "B", "G", "B", "B", "B", "B", "B", "G", "G", 
    "2", "G", "G", "G", "G", "G", "G", "2", "B", "A", "A", "B", "B", "2", 
    "A", "A", "B", "A", "G", "G", "B", "3", "B", "B", "B", "B", "A", "G", 
    "B", "B", "B", "B", "G", "G", "G", "G", "1", "B", "G", "B", "B", "G", 
    "1", "G", "G", "G", "G", "B", "B", "G", "G", "B", "G", "B", "G", "G", 
    "B", "A", "B", "G", "B", "G", "B", "B", "G", "B", "B", "B", "B", "B", 
    "B", "B", "A", "B", "B", "G", "B", "B", "B", "G", "2", "3", "3", "B", 
    "A", "B", "3", "2", "B", "G", "3", "A", "B", "B", "A", "B", "G", "A", 
    "B", "B", "0", "B", "G", "G", "B", "G", "G", "1", "3", "1", "B", "G", 
    "G", "G", "G", "2", "G", "G", "B", "B", "B", "B", "B", "B", "B", "A", 
    "G", "A", "2", "2", "A", "0", "2", "B", "G", "B", "G", "A", "B", "B", 
    "B", "B", "G", "B", "B", "B", "G", "B", "B", "B", "B", "B", "G", "G", 
    "B", "B", "B", "B", "B", "A", "B", "B", "A", "1", "A", "G", "B", "B", 
    "B", "A", "B", "B", "A", "B", "G", "B", "G", "G", "G", "3", "3", "3", 
    "3", "3", "B", "B", "B", "B", "B", "G", "B", "3", "G", "3", "G", "G", 
    "G", "3", "G", "2", "G", "2", "B", "B", "1", "B", "G", "G", "G", "G", 
    "G", "G", "G", "B", "1", "G", "G", "B", "B", "A", "3", "A", "1", "A", 
    "B", "A", "B", "B", "B", "A", "A", "2", "3", "3", "B", "B", "B", "B", 
    "3", "G", "G", "G", "G", "B", "B", "B", "B", "B", "B", "G", "A", "G", 
    "B", "B", "G", "B", "B", "B", "B", "3", "G", "B", "G", "G", "G", "G", 
    "G", "G", "G", "B", "G", "G", "2", "1", "G", "B", "1", "3", "2", "B", 
    "1", "B", "1", "2", "2", "2", "B", "B", "A", "B", "B", "G", "G", "G", 
    "G", "G", "G", "B", "G", "2", "2", "A", "B", "3", "2", "G", "3", "1", 
    "B", "B", "G", "B", "B", "B", "G", "B", "B", "B", "2", "B", "B", "2", 
    "B", "A", "B", "B", "B", "B", "1", "B", "B", "B", "1", "B", "G", "B", 
    "A", "G", "G", "G", "B", "G", "1", "2", "3", "3", "B", "1", "B", "B", 
    "G", "B", "B", "B", "G", "B", "G", "B", "G", "2", "G", "G", "3", "G", 
    "B", "G", "2", "A", "G", "A", "B", "B", "B", "B", "2", "2", "1", "B", 
    "2", "B", "B", "B", "B", "A", "B", "B", "A", "A", "B", "B", "B", "2", 
    "A", "3", "B", "B", "3", "B", "3", "B", "B", "B", "A", "A", "B", "3", 
    "B", "A", "2", "A", "A", "0", "0", "1", "B", "B", "2" ;

 lon = -151.6675, -151.6656, -151.6647, -151.6846, -151.6843, -151.6852, 
    -151.6346, -151.627, -151.5435, -151.5449, -151.5255, -151.5281, 
    -151.5393, -151.5663, -151.5678, -151.5309, -151.5462, -151.5548, 
    -151.5249, -151.5319, -151.5461, -151.5419, -151.5037, -151.5321, 
    -151.5745, -151.5425, -151.538, -151.5453, -151.5504, -151.5424, 
    -151.527, -151.5124, -151.5129, -151.5437, -151.5538, -151.5583, 
    -151.5441, -151.5576, -151.5958, -151.6139, -151.6545, -151.6408, 
    -151.6606, -151.6606, -151.6653, -151.6618, -151.6597, -151.6514, 
    -151.6603, -151.6683, -151.6605, -151.6575, -151.5972, -151.6337, 
    -151.625, -151.6179, -151.6178, -151.6061, -151.5876, -151.5676, 
    -151.5993, -151.5537, -151.5362, -151.6251, -151.5002, -151.487, 
    -151.483, -151.4676, -151.3782, -151.3951, -151.3984, -151.4312, 
    -151.3844, -151.4302, -151.3956, -151.4425, -151.4043, -151.4575, 
    -151.4004, -151.4125, -151.4531, -151.3866, -151.3757, -151.4536, 
    -151.3292, -151.3089, -151.4412, -151.3407, -151.3618, -151.441, 
    -151.3693, -151.4397, -151.3299, -151.3468, -151.3424, -151.3396, 
    -151.3403, -151.344, -151.3497, -151.3564, -151.5106, -151.5712, 
    -151.5787, -151.5812, -151.5851, -151.5989, -151.5378, -151.601, 
    -151.5909, -151.5901, -151.6078, -151.5374, -151.5373, -151.5456, 
    -151.5502, -151.5386, -151.5382, -151.5404, -151.5392, -151.5389, 
    -151.5485, -151.5815, -151.5521, -151.5479, -151.5485, -151.5437, 
    -151.5469, -151.5649, -151.5818, -151.5844, -151.583, -151.5741, 
    -151.5792, -151.5761, -151.5667, -151.546, -151.546, -151.5516, -151.572, 
    -151.5502, -151.5558, -151.5872, -151.5469, -151.5444, -151.5436, 
    -151.5619, -151.6406, -151.5752, -151.5715, -151.5552, -151.5399, 
    -151.5468, -151.5523, -151.5399, -151.5395, -151.5468, -151.5465, 
    -151.543, -151.5341, -151.51, -151.5099, -151.5104, -151.5068, -151.5079, 
    -151.5079, -151.5073, -151.5034, -151.5038, -151.4969, -151.4877, 
    -151.5075, -151.4875, -151.5108, -151.5228, -151.5073, -151.4255, 
    -151.4617, -151.5164, -151.4563, -151.4514, -151.4683, -151.5076, 
    -151.5061, -151.5168, -151.5136, -151.5128, -151.5287, -151.5328, 
    -151.5207, -151.5155, -151.5134, -151.5175, -151.5195, -151.517, 
    -151.5168, -151.5316, -151.5398, -151.5571, -151.5742, -151.5148, 
    -151.6318, -151.6412, -151.6503, -151.6053, -151.6353, -151.6681, 
    -151.6836, -151.6169, -151.6249, -151.6274, -151.6276, -151.6178, 
    -151.6179, -151.6134, -151.5535, -151.5985, -151.5462, -151.563, 
    -151.5729, -151.5565, -151.5534, -151.5694, -151.5876, -151.5855, 
    -151.5721, -151.5722, -151.597, -151.5448, -151.534, -151.5273, 
    -151.3421, -151.3622, -151.1264, -151.1237, -151.1252, -151.1159, 
    -151.1297, -151.1165, -151.1225, -151.1275, -151.1237, -151.1236, 
    -151.1281, -151.1531, -151.1205, -151.1243, -151.1274, -151.1201, 
    -151.123, -151.1235, -151.1072, -151.1058, -151.1048, -151.059, -151.055, 
    -151.5364, -151.5392, -151.5185, -151.5246, -151.531, -151.5085, 
    -151.5105, -151.5229, -151.5247, -151.5353, -151.3849, -151.5284, 
    -151.5314, -151.5294, -151.5462, -151.5782, -151.5661, -151.5945, 
    -151.5954, -151.6044, -151.5961, -151.6353, -151.6297, -151.6647, 
    -151.6576, -151.6894, -151.6609, -151.7119, -151.6609, -151.6586, 
    -151.6505, -151.6498, -151.6605, -151.6664, -151.6516, -151.6662, 
    -151.6712, -151.6472, -151.6768, -151.6373, -151.6424, -151.6338, 
    -151.6294, -151.6777, -151.5549, -151.5412, -151.5286, -151.5152, 
    -151.5061, -151.4941, -151.4989, -151.5046, -151.5207, -151.5092, 
    -151.4925, -151.4884, -151.517, -151.4827, -151.4975, -151.4916, 
    -151.503, -151.5182, -151.5276, -151.5417, -151.7778, -151.5163, 
    -151.4947, -151.4801, -151.4862, -151.4657, -151.5067, -151.5108, 
    -151.5066, -151.5377, -151.5255, -151.4731, -151.475, -151.5013, 
    -151.5014, -151.5101, -151.4933, -151.4706, -151.4875, -151.5089, 
    -151.4922, -151.5154, -151.4892, -151.5083, -151.5198, -151.5079, 
    -151.4873, -151.4992, -151.5031, -151.5235, -151.5343, -151.5471, 
    -151.6552, -151.6605, -151.6525, -151.6501, -151.6532, -151.6446, 
    -151.6622, -151.6641, -151.6647, -151.6638, -151.6655, -151.6646, 
    -151.6635, -151.6556, -151.6608, -151.6607, -151.6633, -151.6594, 
    -151.6583, -151.6463, -151.6516, -151.6599, -151.6614, -151.6628, 
    -151.6579, -151.6564, -151.6488, -151.6401, -151.6454, -151.6379, 
    -151.6307, -151.6311, -151.6288, -151.4243, -151.4274, -151.4279, 
    -151.4521, -151.4495, -151.4813, -151.4998, -151.5235, -151.5301, 
    -151.5084, -151.5135, -151.5198, -151.5269, -151.4782, -151.49, 
    -151.4552, -151.4904, -151.4771, -151.4866, -151.4913, -151.4599, 
    -151.4477, -151.4286, -151.4412, -151.4411, -151.4393, -151.4505, 
    -151.4405, -151.4633, -151.4556, -151.4496, -151.4832, -151.4275, 
    -151.4553, -151.4679, -151.4959, -151.6372, -151.6352, -151.6046, 
    -151.5838, -151.5571, -151.5179, -151.4734, -151.4522, -151.4383, 
    -151.4197, -151.4017, -151.478, -151.4105, -151.3964, -151.3739, 
    -151.4631, -151.3846, -151.3743, -151.3616, -151.3582, -151.3435, 
    -151.3749, -151.3303, -151.2986, -151.3092, -151.2872, -151.2804, 
    -151.2863, -151.2703, -151.2798, -151.3155, -151.3439, -151.3153, 
    -151.3141, -151.3174, -151.3201, -151.2977, -151.3251, -151.4546, 
    -151.3858, -151.3835, -151.3809, -151.513, -151.4372, -151.4416, 
    -151.4491, -151.7043, -151.6881, -151.6641, -151.6509, -151.6424, 
    -151.6407, -151.6408, -151.5081, -151.6411, -151.6319, -151.6004, 
    -151.6538, -151.6646, -151.5791, -151.5687, -151.5654, -151.5675, 
    -151.5675, -151.5706, -151.5958, -151.5052, -151.4841, -151.492, 
    -151.4977, -151.5285, -151.5012, -151.5232, -151.5226, -151.5078, 
    -151.5191, -151.5918, -151.4999, -151.5883, -151.502, -151.5855, 
    -151.5146, -151.5185, -151.5039, -151.5256, -151.5155, -151.4962, 
    -151.4436, -151.5403, -151.5106, -151.5175, -151.4772, -151.4956, 
    -151.4834, -151.4868, -151.4941, -151.4895, -151.4867, -151.4854, 
    -151.4928, -151.4834, -151.4814, -151.4787, -151.4782, -151.4788, 
    -151.4843, -151.4879, -151.4866, -151.4867, -151.4866, -151.4871, 
    -151.4874, -151.488, -151.4884, -151.5042, -151.5357, -151.5602, 
    -151.5892, -151.6291, -151.6526, -151.6607, -151.668, -151.6855, 
    -151.6962, -151.6857, -151.6828, -151.6343, -151.6808, -151.6121, 
    -151.6709, -151.5818, -151.6642, -151.5392, -151.5234, -151.5352, 
    -151.5359, -151.5547, -151.506, -151.5055, -151.5045, -151.49, -151.4875, 
    -151.4945, -151.4868, -151.4878, -151.5019, -151.4931, -151.4866, 
    -151.493, -151.4779, -151.4615, -151.4857, -151.4708, -151.4715, 
    -151.4788, -151.5196, -151.4346, -151.434, -151.4294, -151.4306, 
    -151.4326, -151.4466, -151.4416, -151.4225, -151.4087, -151.3982, 
    -151.4091, -151.5148, -151.7384, -151.6265, -151.5914, -151.5832, 
    -151.5314, -151.5805, -151.5486, -151.5252, -151.5287, -151.5025, 
    -151.4791, -151.5074, -151.5174, -151.5162, -151.5181, -151.5136, 
    -151.5598, -151.562, -151.5955, -151.5747, -151.663, -151.6469, 
    -151.6682, -151.6485, -151.6624, -151.6765, -151.6763, -151.7028, 
    -151.6291, -151.6274, -151.6348, -151.6251, -151.5738, -151.5636, 
    -151.563, -151.5633, -151.5572, -151.5461, -151.4591, -151.3453, 
    -151.3455, -151.3617, -151.3566, -151.307, -151.305, -151.2914, 
    -151.3139, -151.327, -151.3462, -151.2707, -151.2521, -151.3796, 
    -151.3681, -151.365, -151.3643, -151.3602, -151.3781, -151.37, -151.3191, 
    -151.3617, -151.3614, -151.369, -151.378, -151.3713, -151.365, -151.3754, 
    -151.3734, -151.3624, -151.3545, -151.368, -151.3213, -151.3566, 
    -151.3207, -151.3255, -151.3327, -151.2064, -151.2121, -151.2088, 
    -151.2025, -151.2017, -151.2012, -151.2027, -151.2166, -151.2068, 
    -151.2278, -151.2454, -151.2462, -151.2436, -151.2459, -151.2135, 
    -151.2494, -151.2594, -151.2947, -151.3138, -151.3164, -151.3203, 
    -151.3366, -151.338, -151.3594, -151.374, -151.3761, -151.3656, 
    -151.3653, -151.3707, -151.3674, -151.39, -151.3918, -151.3318, 
    -151.3848, -151.2789, -151.299, -151.3016, -151.32, -151.2916, -151.3237, 
    -151.3415, -151.3611, -151.3822, -151.388, -151.434, -151.3685, 
    -151.3808, -151.3615, -151.3778, -151.4126, -151.3705, -151.3625, 
    -151.3623, -151.3621, -151.3568, -151.3664, -151.3586, -151.3623, 
    -151.3604, -151.3605, -151.3628, -151.3902, -151.2628, -151.3701, 
    -151.3745, -151.3482, -151.3683, -151.3614, -151.3589, -151.3588, 
    -151.3672, -151.368, -151.35, -151.3714, -151.3502, -151.3662, -151.3506, 
    -151.3615, -151.3577, -151.362, -151.3592, -151.3646, -151.3539, 
    -151.3563, -151.3731, -151.3608, -151.3607, -151.3649, -151.3609, 
    -151.3614, -151.3765, -151.3971, -151.4391, -151.4533, -151.5005, 
    -151.4659, -151.6037, -151.6334, -151.6487, -151.6621, -151.6569, 
    -151.6382, -151.6585, -151.6263, -151.6342, -151.7576, -151.6586, 
    -151.6422, -151.6624, -151.6628, -151.654, -151.6654, -151.6788, 
    -151.6698, -151.6822, -151.6614, -151.6691, -151.6702, -151.6912, 
    -151.6531, -151.6147, -151.5881, -151.5614, -151.5459, -151.5345, 
    -151.5096, -151.4733, -151.4548, -151.4518, -151.673, -151.5904, 
    -151.3659, -151.3675, -151.3436, -151.3239, -151.2569, -151.3266, 
    -151.3249, -151.2068, -151.2178, -151.1713, -151.1485, -151.1506, 
    -151.1235, -151.1306, -151.1207, -151.111, -151.1131, -151.1137, 
    -151.0834, -151.0809, -151.1118, -150.9977, -151.1111, -151.0918, 
    -151.1197, -151.1871, -151.1897, -151.1633, -151.1676, -151.1814, 
    -151.1812, -151.2113, -151.1894, -151.1904, -151.1902, -151.1913, 
    -151.1974, -151.1908, -151.1488, -151.0803, -151.0817, -151.082, 
    -151.0329, -151.0965, -151.0908, -150.974, -151.0095, -151.1187, 
    -151.1131, -151.0898, -151.0994, -151.1014, -151.1136, -151.1105, 
    -151.107, -151.0618, -151.1968, -151.1963, -151.1673, -151.1855, 
    -151.1799, -151.2333, -151.1794, -151.2372, -151.2372, -151.2371, 
    -151.2455, -151.2539, -151.2546, -151.2488, -151.2493, -151.2497, 
    -151.2439, -151.2448, -151.2748, -151.2885, -151.2201, -151.2305, 
    -151.2352, -151.3223, -151.3426, -151.3486, -151.3613, -151.3503, 
    -151.3595, -151.3659, -151.4216, -151.3761, -151.4378, -151.4189, 
    -151.3966, -151.4387, -151.482, -151.5241, -151.6273, -151.6274, 
    -151.6228, -151.6034, -151.63, -151.6079, -151.5059, -151.4974, 
    -151.3696, -151.3547, -151.2631, -151.1883, -151.194, -151.194, 
    -151.1915, -151.1829, -151.1874, -151.1934, -151.1682, -151.145, 
    -151.1489, -151.1091, -151.1127, -151.1028, -151.1444, -151.1739, 
    -151.1547, -151.2757, -151.3046, -151.328, -151.3415, -151.3531, 
    -151.3595, -151.3516, -151.3345, -151.3189, -151.3001, -151.2786, 
    -151.2044, -151.2119, -151.1366, -151.5456, -151.1967, -151.1946, 
    -151.2084, -151.2007, -151.1991, -151.1977, -151.4999, -151.4989, 
    -151.5187, -151.5069, -151.5129, -151.5218, -151.5109, -151.5139, 
    -151.5008, -151.5059, -151.5146, -151.509, -151.5169, -151.5041, 
    -151.4952, -151.5103, -151.5327, -151.5925, -151.5212, -151.4641, 
    -151.4974, -151.4829, -151.4811, -151.4788, -151.479, -151.4801, 
    -151.4963, -151.508, -151.5228, -151.6224, -151.6405, -151.6414, 
    -151.6604, -151.6625, -151.7092, -151.7086, -151.6617, -151.6764, 
    -151.6703, -151.6591, -151.6582, -151.6667, -151.6667, -151.6735, 
    -151.6585, -151.6583, -151.6583, -151.6589, -151.6647, -151.646, 
    -151.6819, -151.6878, -151.6366, -151.5688, -151.565, -151.5533, 
    -151.5466, -151.5447, -151.5441, -151.5416, -151.5336, -151.5132, 
    -151.5076, -151.5141, -151.499, -151.5091, -151.5202, -151.5255, 
    -151.4921, -151.5314, -151.5284, -151.5224, -151.5108, -151.4924, 
    -151.528, -151.5175, -151.5177, -151.5175, -151.4908, -151.4913, 
    -151.5124, -151.5197, -151.5128, -151.5093, -151.4839, -151.4666, 
    -151.4561, -151.4117, -151.4515, -151.3073, -151.4214, -151.2967, 
    -151.247, -151.4036, -151.3241, -151.3017, -151.3043, -151.1768, 
    -151.2948, -151.1343, -151.1335, -151.1333, -151.0974, -151.1271, 
    -151.1054, -151.0941, -151.0991, -151.0975, -151.0366, -151.0684, 
    -151.0528, -151.0856, -151.0806, -151.0855, -151.0684, -151.076, 
    -151.0999, -150.9906, -151.0957, -151.1286, -151.2186, -151.1859, 
    -151.1861, -151.1885, -151.1601, -151.1589, -151.1791, -151.1869, 
    -151.194, -151.1861, -151.1911, -151.1921, -151.1799, -151.1958, 
    -151.2029, -151.2023, -151.1739, -151.176, -151.1769, -151.1819, 
    -151.1617, -151.1816, -151.1568, -151.1816, -151.2063, -151.1816, 
    -151.1797, -151.1818, -151.185, -151.1531, -151.1286, -151.1472, 
    -151.1624, -151.1903, -151.194, -151.5936, -151.197, -151.2122, 
    -151.2204, -151.2207, -151.2236, -151.2475, -151.2502, -151.2366, 
    -151.2137, -151.2015, -151.2019, -151.202, -151.2015, -151.207, 
    -151.2317, -151.2368, -151.2548, -151.2543, -151.2609, -151.2778, 
    -151.2568, -151.275, -151.3504, -151.3666, -151.4765, -151.4985, 
    -151.545, -151.5, -151.5364, -151.5311, -151.551, -151.5502, -151.5526, 
    -151.5167, -151.5124, -151.5024, -151.485, -151.4877, -151.4917, 
    -151.4949, -151.4868, -151.4999, -151.4946, -151.4943, -151.5111, 
    -151.5044, -151.4948, -151.4948, -151.4991, -151.4931, -151.4927, 
    -151.4946, -151.4962, -151.4958, -151.4973, -151.5113, -151.4967, 
    -151.487, -151.502, -151.5034, -151.5181, -151.5012, -151.5355, -151.5, 
    -151.5051, -151.5445, -151.5765, -151.5793, -151.2171, -151.2017, 
    -151.2021, -151.202, -151.252, -151.2889, -151.3002, -151.6397, 
    -151.5662, -151.5368, -151.2382, -151.2325, -151.1974, -151.1724, 
    -151.1869, -151.186, -151.182, -151.1825, -151.1746, -151.1873, 
    -151.1699, -151.192, -151.1883, -151.1991, -151.1865, -151.1841, 
    -151.1817, -151.1855, -151.2017, -151.2196, -151.2123, -151.2166, 
    -151.2132, -151.2159, -151.2109, -151.2158, -151.3863, -151.4283, 
    -151.1996, -151.5133, -151.5291, -151.2587, -151.2709, -151.5296, 
    -151.5792, -151.6394, -151.5832, -151.9322, -151.6305, -151.5774, 
    -151.5989, -151.708, -151.5696, -151.739, -151.5726, -151.6216, 
    -151.5851, -151.5666, -151.5863, -151.6693, -151.9277, -151.6656, 
    -151.6406, -151.6396, -151.6568, -151.6482, -151.6877, -151.6616, 
    -151.6044, -151.6625, -151.6708, -151.7043, -151.6546, -151.6543, 
    -151.6485, -151.6704, -151.6684, -151.669, -151.6826, -151.6628, 
    -151.6493, -151.6736, -151.6325, -151.6366, -151.6261, -151.6544, 
    -151.6147, -151.5666, -151.5663, -151.5662, -151.566, -151.5658, 
    -151.5276, -151.586, -151.5856, -151.58, -151.5802, -151.5786, -151.5512, 
    -151.5742, -151.5688, -151.6017, -151.5626, -151.533, -151.5682, 
    -151.5689, -151.5577, -151.5779, -151.569, -151.5699, -151.5766, 
    -151.579, -151.5738, -151.5764, -151.576, -151.5668, -151.5688, 
    -151.5706, -151.5753, -151.5683, -151.5815, -151.5719, -151.5812, 
    -151.5667, -151.5928, -151.57, -151.5755, -151.5685, -151.5663, 
    -151.5386, -151.6173, -151.5384, -151.5368, -151.5775, -151.6014, 
    -151.6338, -151.6393, -151.6795, -151.6615, -151.6673, -151.6576, 
    -151.6692, -151.6654, -151.661, -151.6707, -151.6893, -151.6797, 
    -151.6604, -151.6507, -151.6502, -151.6684, -151.6455, -151.656, 
    -151.6645, -151.6749, -151.6619, -151.6588, -151.6063, -151.4796, 
    -151.5295, -151.531, -151.487, -151.5268, -151.5305, -151.5017, 
    -151.5342, -151.5257, -151.5352, -151.5169, -151.5393, -151.5178, 
    -151.5387, -151.5242, -151.5084, -151.4987, -151.5004, -151.4529, 
    -151.459, -151.4595, -151.4604, -151.4692, -151.4693, -151.3881, 
    -151.4807, -151.4927, -151.4806, -151.4706, -151.4762, -151.4609, 
    -151.4573, -151.4468, -151.4614, -151.4429, -151.4319, -151.4427, 
    -151.4333, -151.4468, -151.4572, -151.4697, -151.4456, -151.4702, 
    -151.4681, -151.409, -151.4051, -151.3985, -151.3945, -151.3675, 
    -151.3504, -151.3645, -151.369, -151.3621, -151.3812, -151.3619, 
    -151.406, -151.3719, -151.4294, -151.3637, -151.4489, -151.4696, 
    -151.4861, -151.5173, -151.5369, -151.3607, -151.5569, -151.5363, 
    -151.5713, -151.6768, -151.6902, -151.6951, -151.6896, -151.691, 
    -151.6681, -151.6357, -151.6301, -151.6508, -151.6583, -151.6549, 
    -151.6645, -151.6587, -151.6628, -151.5882, -151.6236, -151.64, 
    -151.6623, -151.6436, -151.6231, -151.652, -151.6709, -151.6702, 
    -151.6574, -151.67, -151.6752, -151.6586, -151.6831, -151.6841, 
    -151.6745, -151.6746, -151.6594, -151.6593, -151.645, -151.6487, 
    -151.6747, -151.6811, -151.6244, -151.6176, -151.4533, -151.369, 
    -151.4142, -151.392, -151.3908, -151.3906, -151.3868, -151.3734, 
    -151.3643, -151.3632, -151.357, -151.4066, -151.3397, -151.3542, 
    -151.3827, -151.438, -151.4402, -151.4268, -151.4355, -151.4355, 
    -151.3941, -151.3903, -151.3338, -151.3609, -151.3688, -151.3644, 
    -151.3663, -151.3647, -151.289, -151.3262, -151.3105, -151.3006, 
    -151.3235, -151.2885, -151.2641, -151.2911, -151.2919, -151.2853, 
    -151.1878, -151.1871, -151.282, -151.2464, -151.0986, -151.1133, 
    -151.0856, -151.1239, -151.1239, -151.1941, -151.1638, -151.2215, 
    -151.1776, -151.1721, -151.1868, -151.4068, -151.4045, -151.4025, 
    -151.3765, -151.3712, -151.5367, -151.4174, -151.4471, -151.4523, 
    -151.4711, -151.4418, -151.4288, -151.4292, -151.4079, -151.4237, 
    -151.4254, -151.3846, -151.3887, -151.3902, -151.4407, -151.3933, 
    -151.4835, -151.482, -151.4746, -151.4981, -151.4997, -151.4664, 
    -151.4697, -151.4717, -151.5321, -151.5206, -151.5028, -151.4875, 
    -151.4959, -151.4681, -151.4874, -151.5224, -151.488, -151.4516, 
    -151.5421, -151.5674, -151.578, -151.5805, -151.5892, -151.57, -151.5367, 
    -151.4902, -151.523, -151.4998, -151.5215, -151.5207, -151.4955, 
    -151.4957, -151.4975, -151.495, -151.4931, -151.3849, -151.39, -151.4423, 
    -151.432, -151.4302, -151.4133, -151.4328, -151.4075, -151.4209, 
    -151.4483, -151.64, -151.6587, -151.6602, -151.6602, -151.66, -151.6599, 
    -151.6592, -151.6513, -151.6614, -151.6252, -151.6599, -151.5981, 
    -151.662, -151.6627, -151.6554, -151.6689, -151.6632, -151.6683, 
    -151.6609, -151.6567, -151.6549, -151.6638, -151.6646, -151.6583, 
    -151.6676, -151.6617, -151.6617, -151.6603, -151.6642, -151.6352, 
    -151.6153, -151.6521, -151.6564, -151.6874, -151.6857, -150.9142, 
    -151.2908, -151.0384, -150.9982, -150.993, -150.9708, -151.1395, 
    -151.0283, -151.0249, -151.0263, -151.0179, -151.0121, -151.0142, 
    -150.9468, -151.0153, -151.022, -151.0158, -151.0206, -151.0131, 
    -151.0137, -150.9922, -151.0135, -151.0151, -151.0433, -151.0397, 
    -151.1257, -151.13, -151.1586, -151.1868, -151.2169, -151.2422, 
    -151.2726, -151.2951, -151.3044, -151.3147, -151.4241, -151.4413, 
    -151.4414, -151.36, -151.4408, -151.449, -151.4482, -151.4408, -151.4338, 
    -151.4703, -151.4936, -151.4739, -151.4853, -151.4707, -151.4584, 
    -151.4413, -151.4562, -151.4501, -151.4501, -151.4451, -151.4472, 
    -151.4603, -151.4602, -151.4467, -151.4568, -151.4403, -151.4424, 
    -151.4405, -151.4622, -151.4551, -151.4394, -151.4481, -151.4532, 
    -151.4697, -151.4415, -151.4431, -151.4427, -151.5264, -151.4879, 
    -151.5056, -151.4859, -151.4221, -151.4029, -151.4228, -151.4328, 
    -151.4101, -151.4264, -151.4284, -151.4321, -151.5365, -151.5513, 
    -151.5745, -151.7255, -151.7281, -151.7468, -151.645, -151.645, 
    -151.6349, -151.6487, -151.6622, -151.6575, -151.6531, -151.6631, 
    -151.6594, -151.6461, -151.6558, -151.6682, -151.6634, -151.6591, 
    -151.6637, -151.6533, -151.6729, -151.6782, -151.651, -151.6586, 
    -151.3898, -151.5559, -151.5893, -151.5995, -151.6328, -151.6445, 
    -151.6194, -151.6619, -151.6601, -151.613, -151.6567, -151.6471, 
    -151.6459, -151.6468, -151.651, -151.6485, -151.6496, -151.6756, 
    -151.6688, -151.6613, -151.6749, -151.661, -151.6732, -151.6657, 
    -151.6664, -151.6702, -151.6439, -151.66, -151.6613, -151.6671, 
    -151.6556, -151.6522, -151.6575, -151.6579, -151.6648, -151.5778, 
    -151.5712, -151.5315, -151.5242, -151.513, -151.3966, -151.3563, 
    -151.3034, -151.283, -151.2877, -151.4654, -151.3022, -151.3022, 
    -151.3197, -151.3127, -151.3191, -151.2842, -151.3087, -151.2987, 
    -151.3116, -151.3248, -151.2991, -151.3147, -151.3051, -151.3106, 
    -151.281, -151.3187, -151.2616, -151.3119, -151.2679, -151.229, 
    -151.2297, -151.2205, -151.2079, -151.1215, -151.1117, -151.1173, 
    -151.117, -151.1173, -151.1188, -151.131, -151.152, -151.3692, -151.3577, 
    -151.3439, -151.3209, -151.3244, -151.3604, -151.3727, -151.3573, 
    -151.3599, -151.3535, -151.3515, -151.3092, -151.3088, -151.2359, 
    -151.2003, -151.2222, -151.2452, -151.2377, -151.223, -151.2185, 
    -151.229, -151.2284, -151.2524, -151.2368, -151.2475, -151.2471, 
    -151.2477, -151.2518, -151.2445, -151.245, -151.2347, -151.2315, 
    -151.2214, -151.1991, -150.9784, -150.9669, -150.9688, -150.9662, 
    -150.9385, -150.9509, -150.9426, -150.9562, -150.9487, -150.9477, 
    -150.9458, -150.9805, -150.9463, -150.982, -150.9773, -150.9809, 
    -150.9821, -150.9071, -150.929, -150.9254, -150.9849, -150.9814, 
    -151.1692, -151.3861, -151.4253, -151.5357, -151.5368, -151.5432, 
    -151.5437, -151.6051, -151.6643, -151.6584, -151.6615, -151.6606, 
    -151.6605, -151.6578, -151.6546, -151.6711, -151.6595, -151.6567, 
    -151.6587, -151.66, -151.6599, -151.6728, -151.6367, -151.6472, 
    -151.6816, -151.6898, -151.7073, -151.7226, -151.7353, -151.6856, 
    -151.6602, -151.6166, -151.6305, -151.6491, -151.6239, -151.6562, 
    -151.667, -151.675, -151.6863, -151.6687, -151.6731, -151.7397, 
    -151.7542, -151.735, -151.74, -151.7659, -151.7289, -151.7544, -151.7462, 
    -151.6635, -151.6718, -151.6793, -151.6725, -151.6605, -151.6606, 
    -151.7188, -151.6703, -151.6665, -151.6417, -151.6372, -151.6537, 
    -151.6571, -151.6574, -151.6626, -151.6001, -151.6165, -151.6156, 
    -151.6108, -151.6001, -151.5717, -151.515, -151.5102, -151.4471, 
    -151.4807, -151.4653, -151.4498, -151.2844, -151.2845, -151.2573, 
    -151.2227, -151.1366, -151.0311, -151.1182, -151.0146, -151.0025, 
    -151.0283, -150.952, -150.9538, -151.0164, -150.8978, -150.9839, -151.06, 
    -151.0485, -151.0437, -151.0358, -151.0119, -151.04, -151.0267, 
    -151.0176, -151.0179, -150.9691, -150.9647, -150.967, -150.9517, 
    -150.9666, -150.9258, -150.9662, -150.943, -150.9636, -151.0208, 
    -150.9578, -151.017, -150.9865, -150.9561, -150.9535, -150.9791, 
    -150.9785, -150.9628, -150.9347, -150.9137, -150.909, -150.91, -150.9262, 
    -150.9081, -150.8861, -150.9071, -150.9066, -150.8986, -150.9113, 
    -150.9125, -150.9035, -150.9193, -150.9157, -150.9267, -150.9227, 
    -150.9154, -150.8938, -150.919, -150.9189, -150.9193, -150.9198, 
    -150.9197, -150.9228, -150.9315, -150.8994, -150.9164, -150.9076, 
    -150.9126, -150.9119, -150.9286, -150.9295, -150.8486, -150.8948, 
    -150.9129, -150.9101, -150.9105, -150.9057, -150.9033, -150.8835, 
    -150.8997, -150.9169, -150.918, -150.9246, -150.9159, -150.9216, 
    -150.9235, -150.9147, -150.9132, -150.9118, -150.9179, -150.9127, 
    -150.9035, -150.9056, -150.9079, -150.9185, -150.9185, -150.9075, 
    -150.8539, -150.8451, -150.9077, -150.9169, -150.9099, -150.9097, 
    -150.9089, -150.9115, -150.9127, -150.9213, -150.9216, -150.9211, 
    -150.9267, -150.9499, -150.9491, -150.9372, -150.9453, -150.9196, 
    -150.9314, -150.9273, -150.9165, -150.9167, -150.9046, -150.9103, 
    -150.9058, -150.9124, -150.9087, -150.9196, -150.9198, -150.9362, 
    -150.9091, -150.9486, -150.909, -150.9491, -150.8922, -150.8922, 
    -150.8983, -150.9004, -150.8978, -150.8868, -150.8882, -150.8754, 
    -150.8762, -150.8459, -150.9193, -150.872, -150.9149, -150.9162, 
    -150.9176, -150.9316, -150.9192, -150.9145, -150.9117, -150.9639, 
    -150.9162, -150.9226, -150.9196, -150.9135, -150.912, -150.904, 
    -150.9032, -150.9183, -150.9046, -150.9032, -150.8621, -150.9155, 
    -150.8929, -150.9115, -150.9043, -150.906, -150.9119, -150.9045, 
    -150.9267, -150.9285, -150.8935, -150.9274, -150.9279, -150.9319, 
    -150.9181, -150.9155, -150.9181, -150.9255, -150.9151, -150.9269, 
    -150.9262, -150.9252, -150.934, -150.9338, -150.9341, -150.9476, 
    -150.9461, -150.9399, -150.8997, -150.9088, -150.9415, -150.9189, 
    -150.9299, -150.9443, -150.9128, -150.9454, -150.9457, -150.9441, 
    -150.9185, -150.95, -150.9578, -151.1798, -151.2716, -151.2463, 
    -151.1582, -151.0541, -151.0583, -151.0418, -150.9952, -151.0305, 
    -150.9641, -150.9322, -150.9208, -150.945, -150.9411, -150.941, 
    -150.8986, -150.9404, -150.8974, -150.9528, -150.9377, -150.9353, 
    -150.9194, -150.8769, -150.8948, -150.927, -150.9243, -150.9249, 
    -150.9301, -150.9269, -150.9638, -150.9274, -150.9376, -150.9397, 
    -150.941, -150.9303, -150.9127, -150.9358, -150.9129, -150.9375, 
    -150.9171, -150.9176, -150.9178, -150.9241, -150.9156, -150.9066, 
    -150.9053, -150.9034, -150.9053, -150.9067, -151.0186, -150.9733, 
    -150.9645, -150.9103, -150.9213, -150.8831, -150.873, -150.8765, 
    -150.9207, -150.9072, -150.8827, -150.8849, -150.9242, -150.9134, 
    -150.8921, -150.8978, -150.9117, -150.9098, -150.881, -150.909, 
    -150.9151, -150.8909, -150.8925, -150.8833, -150.9108, -150.8825, 
    -150.8318, -150.8573, -150.8754, -151.4414, -151.4565, -151.4736, 
    -151.5415, -151.5488, -151.5499, -151.5458, -151.6481, -151.6161, 
    -151.65, -151.6458, -151.6511, -151.6598, -151.6564, -151.6871, 
    -151.6639, -151.6756, -151.6606, -151.6605, -151.698, -151.6629, 
    -151.6601, -151.5358, -151.5774, -151.5663, -151.6545, -151.6443, 
    -151.6615, -151.6608, -151.6642, -151.6637, -151.6498, -151.6583, 
    -151.66, -151.6763, -151.6773, -151.7052, -151.6674, -151.6763, 
    -151.7448, -151.6712, -151.6437, -151.6507, -151.6674, -151.6637, 
    -151.6483, -151.6502, -151.651, -151.7004, -151.6625, -151.6978, 
    -151.661, -151.6564, -151.654, -151.6054, -151.5694, -151.5607, 
    -151.5408, -151.5156, -151.489, -151.4647, -151.4423, -151.612, 
    -151.3797, -151.3075, -151.31, -151.0327, -150.9986, -150.9811, 
    -150.9417, -150.8954, -150.9198, -150.8475, -150.7642, -150.8491, 
    -150.9392, -150.9501, -150.9626, -150.9424, -150.9099, -150.9722, 
    -150.967, -150.9285, -150.956, -150.9493, -150.9185, -150.9612, 
    -151.0404, -151.0142, -151.0391, -151.037, -151.037, -151.0409, 
    -151.0185, -151.052, -151.0594, -151.0642, -151.0096, -151.0489, 
    -151.0894, -151.0856, -151.056, -151.124, -151.0586, -151.058, -151.1459, 
    -151.2203, -151.3455, -151.3623, -151.378, -151.3991, -151.3976, 
    -151.3796, -151.3262, -151.3293, -151.3284, -151.3261, -151.3287, 
    -151.3861, -151.315, -151.3163, -151.3219, -151.4086, -151.4115, 
    -151.3992, -151.3934, -151.455, -151.4538, -151.4372, -151.4477, 
    -151.4451, -151.4425, -151.4426, -151.4441, -151.4414, -151.4517, 
    -151.4429, -151.4398, -151.4608, -151.4101, -151.3594, -151.3164, 
    -151.3188, -151.4008, -151.3171, -151.3877, -151.317, -151.3508, 
    -151.3477, -151.3678, -151.369, -151.3768, -151.3504, -151.3548, 
    -151.3787, -151.382, -151.3603, -151.3607, -151.3469, -151.3608, 
    -151.3988, -151.3828, -151.3889, -151.3981, -151.3993, -151.3892, 
    -151.3891, -151.3979, -151.3889, -151.3878, -151.3876, -151.388, 
    -151.3866, -151.3907, -151.4355, -151.4193, -151.4378, -151.3902, 
    -151.3957, -151.3983, -151.3682, -151.3672, -151.3672, -151.3293, 
    -151.3485, -151.3469, -151.3438, -151.334, -151.2754, -151.2469, 
    -151.2543, -151.2486, -151.2224, -151.2495, -151.2273, -151.2189, 
    -151.2465, -151.2494, -151.1804, -151.245, -151.246, -151.1625, 
    -151.1478, -151.113, -151.2379, -151.231, -151.24, -151.0094, -150.9785, 
    -151.0555, -151.2258, -151.2696, -151.2877, -151.2986, -151.364, 
    -151.1767, -151.1302, -151.4535, -151.4608, -151.4694, -151.4668, 
    -151.4681, -151.4722, -151.4765, -151.4645, -151.4866, -151.4759, 
    -151.5789, -151.6648, -151.5674, -151.5384, -151.5609, -151.5949, 
    -151.5825, -151.6318, -151.6626, -151.6658, -151.6567, -151.6567, 
    -151.7288, -151.6598, -151.6614, -151.6608, -151.6648, -151.5814, 
    -151.6693, -151.7893, -151.6619, -151.6625, -151.6716, -151.6575, 
    -151.6622, -151.6617, -151.6639, -151.6602, -151.662, -151.6605, 
    -151.6649, -151.6876, -151.6672, -151.6617, -151.6693, -151.6621, 
    -151.7029, -151.6824, -151.6555, -151.661, -151.6491, -151.6231, 
    -151.6429, -151.639, -151.639, -151.7102, -151.6025, -151.5972, -151.598, 
    -151.5665, -151.5619, -151.567, -151.5665, -151.5508, -151.4575, 
    -151.3996, -151.41, -151.4062, -151.3093, -151.4445, -151.3438, 
    -151.3296, -151.2996, -151.4329, -151.424, -151.2119, -151.2112, 
    -151.2021, -151.2047, -151.1861, -151.2103, -151.1721, -151.175, 
    -151.2596, -151.2213, -151.2091, -151.1669, -151.1864, -151.2081, 
    -151.2105, -151.1702, -151.1868, -151.1792, -151.1631, -151.1681, 
    -151.1729, -151.1866, -151.1833, -151.1954, -151.191, -151.1874, 
    -151.189, -151.1866, -151.1866, -151.1856, -151.1871, -151.1696, 
    -151.147, -151.1059, -151.161, -151.1613, -151.0244, -151.0257, 
    -151.0194, -151.1525, -151.0159, -151.0343, -151.1275, -150.9758, 
    -151.0155, -151.0214, -151.023, -151.0233, -151.0573, -151.0124, 
    -151.0375, -151.0248, -150.9879, -151.023, -150.9958, -150.9797, 
    -151.0091, -150.9595, -151.0251, -151.0161, -150.9368, -151.0058, 
    -150.9978, -150.9954, -150.9637, -150.9698, -150.9824, -150.9736, 
    -150.9437, -150.9873, -150.9925, -150.9917, -151.0004, -151.0199, 
    -151.0225, -151.0195, -150.948, -151.0158, -150.8924, -151.0158, 
    -151.0333, -151.032, -151.0158, -151.0328, -151.0304, -151.0074, 
    -151.0129, -151.0269, -151.0164, -151.0171, -151.0159, -150.9844, 
    -151.0033, -151.0031, -151.0186, -150.9725, -150.9678, -151.0305, 
    -150.9907, -151.0054, -151.0193, -151.0149, -151.0105, -151.015, 
    -151.0093, -151.0147, -151.022, -151.0263, -151.0322, -151.0268, 
    -151.0373, -151.025, -150.9403, -151.0146, -151.0193, -150.9793, 
    -150.9721, -150.965, -150.9628, -150.961, -150.9768, -150.9641, 
    -150.9627, -150.9547, -150.9658, -150.9667, -150.9697, -150.9803, 
    -150.9751, -150.9752, -150.9727, -150.9688, -150.9591, -150.9573, 
    -150.9799, -150.9892, -150.9738, -150.973, -150.9769, -150.9901, 
    -150.9779, -150.9375, -150.97, -150.9665, -150.9714, -150.9715, 
    -150.9704, -150.9705, -150.972, -150.971, -150.9772, -150.9852, 
    -150.9822, -150.9742, -150.9683, -150.9677, -151.0025, -150.9717, 
    -150.9747, -150.9605, -150.9716, -150.9729, -150.9565, -150.9651, 
    -150.9632, -150.9796, -150.966, -150.9816, -150.9899, -150.9895, 
    -150.9717, -150.9719, -150.9661, -150.9673, -150.9661, -150.9722, 
    -150.9729, -150.9776, -150.9795, -150.9764, -150.9747, -151.0731, 
    -151.08, -151.097, -151.0188, -151.1134, -151.1575, -151.2279, -151.2319, 
    -151.2302, -151.2556, -151.2872, -151.2726, -151.2695, -151.2731, 
    -151.2721, -151.3267, -151.3562, -151.3877, -151.3378, -151.3585, 
    -151.3511, -151.3698, -151.4213, -151.4677, -151.4849, -151.489, 
    -151.5084, -151.5554, -151.6497, -151.6548, -151.6712, -151.9516, 
    -151.6603, -151.6449, -151.6649, -151.656, -151.6656, -151.6555, 
    -151.6628, -151.6651, -151.6676, -151.6436, -151.6437, -151.6574, 
    -151.6608, -151.6505, -151.6499, -151.6552, -151.6812, -151.7074, 
    -151.6442, -151.6339, -151.6038, -151.6294, -151.2221, -151.1453, 
    -151.1972, -151.2147, -151.4203, -151.4422, -151.4587, -151.481, 
    -151.6281, -151.6458, -151.6588, -151.6347, -151.6559, -151.6567, 
    -151.6776, -151.6786, -151.6244, -151.6617, -151.6227, -151.6926, 
    -151.719, -151.7214, -151.717, -151.6891, -151.7021, -151.7198, 
    -151.7012, -151.6917, -151.7163, -151.7065, -151.6992, -151.7114, 
    -151.6988, -151.6935, -151.6945, -151.701, -151.6963, -151.6966, 
    -151.6965, -151.6396, -151.7301, -151.7613, -151.6933, -151.5412, 
    -151.4143, -151.6101, -151.6795, -151.375, -151.3665, -151.6946, 
    -151.3455, -151.3355, -151.6713, -151.591, -151.5891, -151.2623, 
    -151.2758, -151.2681, -151.2484, -151.2288, -151.2607, -151.2383, 
    -151.2309, -151.2384, -151.2356, -151.2382, -151.2462, -151.2401, 
    -151.242, -151.2424, -151.2456, -151.2236, -151.1813, -151.1888, 
    -151.1859, -151.1852, -151.1271, -150.9627, -150.9658, -150.9632, 
    -150.9636, -150.9638, -150.9641, -150.8275, -151.0126, -151.024, 
    -151.0235, -150.9952, -150.9939, -150.9992, -151.0079, -151.0152, 
    -151.0211, -151.0143, -151.0151, -151.0072, -151.0069, -151.017, 
    -151.031, -151.0191, -151.0303, -151.0179, -151.029, -151.0174, -151.029, 
    -151.1317, -151.0507, -151.018, -151.0566, -151.0547, -151.0508, 
    -151.0509, -151.0511, -151.0508, -151.0281, -151.0298, -151.0334, 
    -151.0318, -151.0312, -151.0418, -151.0124, -151.0385, -151.0365, 
    -151.0436, -151.0123, -151.0169, -151.067, -151.013, -150.9736, 
    -150.9642, -150.95, -150.9865, -150.9607, -150.9738, -150.9917, 
    -150.9991, -150.9952, -150.9974, -150.9957, -150.9648, -150.969, 
    -150.9686, -150.9686, -150.9689, -150.9689, -150.9688, -150.9902, 
    -150.9931, -150.9693, -150.9694, -150.9674, -150.9694, -150.9529, 
    -151.0051, -151.006, -150.9913, -151.0215, -151.026, -151.0282, -151.026, 
    -151.0306, -151.0055, -151.0178, -151.0062, -151.0171, -151.0114, 
    -151.0208, -150.9738, -150.9347, -150.9326, -150.972, -150.9215, 
    -151.0084, -151.3893, -151.4568, -151.4652, -151.4809, -151.4066, 
    -151.6614, -151.7019, -151.673, -151.6495, -151.6513, -151.6548, 
    -151.6575, -151.6692, -151.6568, -151.6602, -151.6562, -151.6545, 
    -151.6519, -151.6626, -151.6624, -151.6612, -151.659, -151.6589, 
    -151.6608, -151.662, -151.6737, -151.6777, -151.212, -151.2109, 
    -151.2162, -151.2126, -151.1965, -151.1554, -151.1934, -151.1867, 
    -151.1871, -151.1821, -151.1612, -151.1514, -151.1304, -151.1194, 
    -151.2022, -151.1169, -151.1085, -151.1291, -151.0779, -151.0633, 
    -151.0528, -151.0472, -151.0487, -151.0296, -150.9997, -151.0273, 
    -150.986, -150.9962, -150.9964, -151.0139, -151.0135, -150.9815, 
    -150.9679, -150.9915, -150.9985, -150.9887, -151.0252, -150.9837, 
    -150.9682, -150.9709, -150.9605, -150.979, -150.9497, -150.9666, 
    -150.963, -150.9626, -150.9655, -150.9667, -150.9675, -150.9736, 
    -150.966, -151.0584, -150.9785, -151.0553, -151.0646, -151.0571, 
    -150.9687, -150.976, -151.0225, -151.0188, -151.0363, -151.0796, 
    -151.0584, -151.1303, -151.1133, -151.0943, -151.0914, -151.1021, 
    -151.118, -151.1628, -151.1741, -151.206, -151.1876, -151.257, -151.255, 
    -151.2497, -150.924, -151.2644, -151.2459, -151.2345, -151.2568, 
    -151.2618, -151.2579, -151.2586, -151.2574, -151.2451, -151.2588, 
    -151.2558, -151.2574, -151.2609, -151.2602, -151.259, -151.2231, 
    -151.1971, -151.2207, -151.2036, -151.1984, -151.1869, -151.1749, 
    -151.1355, -151.1323, -151.1152, -151.118, -151.0918, -151.0729, 
    -151.0736, -151.0736, -151.0655, -150.9925, -151.1751, -150.967, 
    -151.2229, -151.2151, -151.2081, -151.2147, -151.2155, -151.2245, 
    -151.2313, -151.2583, -151.3545, -151.3585, -151.3426, -151.3283, 
    -151.3082, -151.2939, -151.3004, -151.3104, -151.2648, -151.4431, 
    -151.3581, -151.3484, -151.3481, -151.3452, -151.3648, -151.365, 
    -151.3671, -151.3658, -151.3813, -151.3998, -151.3593, -151.4238, 
    -151.4402, -151.4667, -151.4854, -151.4503, -151.4993, -151.5162, 
    -151.4971, -151.5285, -151.549, -151.5835, -151.5806, -151.6385, 
    -151.5792, -151.5825, -151.5741, -151.5831, -151.6452, -151.6389, 
    -151.6393, -151.6747, -151.6873, -151.5483, -151.557, -151.4343, 
    -151.3933, -151.3955, -151.3529, -151.3522, -151.3492, -151.3206, 
    -151.3138, -151.2893, -151.3157, -151.3165, -151.2512, -151.2661, 
    -151.3193, -151.2883, -151.2698, -151.2713, -151.2306, -151.2493, 
    -151.2387, -151.2375, -151.2068, -151.1626, -151.1854, -151.1854, 
    -151.1035, -151.2874, -151.1959, -151.1967, -151.2432, -151.2451, 
    -151.1773, -151.165, -151.1326, -151.2083, -151.1998, -151.2093, 
    -151.1041, -151.0913, -151.0909, -151.0976, -151.0916, -151.0539, 
    -151.0549, -151.033, -151.0341, -151.029, -151.0282, -151.0273, 
    -151.0099, -151.0127, -151.0125, -151.0087, -151.0236, -150.9453, 
    -150.9451, -151.0106, -151.0105, -151.0012, -151.0152, -151.0255, 
    -151.091, -151.1057, -151.3655, -151.3832, -151.4091, -151.413, 
    -151.2133, -151.2223, -151.4007, -151.3005, -151.3972, -151.4065, 
    -151.4134, -151.2921, -151.3114, -151.3064, -151.3129, -151.3765, 
    -151.332, -151.328, -151.3234, -151.3159, -151.3025, -151.2995, 
    -151.2633, -151.2258, -151.1886, -151.1902, -151.1805, -151.1658, 
    -151.1684, -151.1427, -151.1326, -151.1595, -151.1199, -151.0419, 
    -151.016, -151.0151, -150.975, -150.9743, -151.0311, -151.0802, 
    -150.9577, -151.1368, -151.1265, -151.1867, -151.1537, -151.1909, 
    -151.2329, -151.6381, -151.6378, -151.6356, -151.6398, -151.6644, 
    -151.649, -151.6584, -151.6988, -151.6436, -151.6671, -151.6724, 
    -151.6767, -151.6636, -151.6373, -151.644, -151.6469, -151.6548, 
    -151.6515, -151.6573, -151.6593, -151.6563, -151.675, -151.6899, 
    -151.7006, -151.7119, -151.7173, -151.8129, -151.8607, -151.6396, 
    -151.6455, -151.8782, -151.8705, -151.8645, -151.8283, -151.8599, 
    -151.8282, -151.9151, -151.791, -151.7882, -151.7758, -151.7729, 
    -151.8132, -151.7749, -151.7775, -151.8007, -151.7537, -151.7468, 
    -151.7516, -151.7628, -151.774, -151.7759, -151.7427, -151.7037, 
    -151.7157, -151.708, -151.7143, -151.7138, -151.7109, -151.6859, 
    -151.661, -151.6527, -151.6433, -151.6299, -151.6119, -151.5503, 
    -151.5927, -151.398, -151.3852, -151.351, -151.3383, -151.3382, 
    -151.3431, -151.321, -151.309, -151.2987, -151.2488, -151.2189, 
    -151.2078, -151.1969, -151.1967, -151.155, -151.458, -151.4616, 
    -150.9992, -150.9964, -151.0191, -150.9902, -150.995, -150.9872, 
    -150.9836, -150.9781, -150.9778, -150.9324, -150.9575, -150.9421, 
    -150.9438, -150.9438, -150.971, -151.0607, -151.0368, -151.0853, 
    -151.1297, -150.9712, -151.0995, -150.9288, -150.9471, -151.0749, 
    -151.0141, -151.0213, -150.9917, -151.0027, -150.9847, -150.9717, 
    -150.9732, -150.97, -150.9574, -150.9484, -150.9652, -150.9589, 
    -150.9563, -150.9604, -150.9601, -150.9601, -150.9621, -150.9654, 
    -150.9617, -150.9653, -150.9647, -150.9693, -150.9653, -150.9645, 
    -150.9686, -150.9695, -150.976, -150.983, -150.981, -150.9744, -150.9667, 
    -150.9655, -150.965, -150.965, -150.9649, -150.9661, -150.9681, 
    -150.9688, -150.9712, -150.9733, -150.975, -150.9778, -150.9826, 
    -150.9874, -150.9865, -150.9869, -151.003, -151.0058, -151.0099, 
    -151.0122, -151.0125, -151.0107, -151.0082, -151.0131, -151.0075, 
    -151.0347, -151.0432, -151.0233, -151.0356, -151.0267, -151.0362, 
    -151.1044, -151.1887, -151.178, -151.2208, -151.299, -151.3218, 
    -151.3419, -151.3986, -151.3849, -151.404, -151.4076, -151.4262, 
    -151.4357, -151.4367, -151.4465, -151.4431, -151.4472, -151.4621, 
    -151.4406, -151.4384, -151.4447, -151.4511, -151.477, -151.4607, 
    -151.4581, -151.4635, -151.4679, -151.479, -151.4949, -151.4776, 
    -151.5124, -151.5174, -151.5228, -151.5427, -151.5592, -151.5313, 
    -151.5649, -151.6336, -151.593, -151.6356, -151.6218, -151.6611, 
    -151.6605, -151.661, -151.6589, -151.6616, -151.9827, -151.6741, 
    -151.6575, -151.6534, -151.6598, -151.6621, -151.6611, -151.6571, 
    -151.6522, -151.667, -151.6635, -151.6675, -151.661, -151.6639, 
    -151.7446, -151.642, -151.6381, -151.6275, -151.6283, -151.6319, 
    -151.6758, -151.6355, -151.6339, -151.6271, -151.6193, -151.6004, 
    -151.541, -151.5425, -151.5452, -151.5442, -151.5456, -151.5156, 
    -151.4916, -151.5391, -151.4762, -151.5371, -151.584, -151.4587, 
    -151.582, -151.518, -151.4358, -151.4093, -151.4329, -151.3819, 
    -151.4297, -151.3845, -151.3364, -151.3256, -151.3255, -151.2937, 
    -151.2956, -151.2379, -151.2569, -151.2542, -151.264, -151.269, 
    -151.2569, -151.2637, -151.2577, -151.2386, -151.2476, -151.2461, 
    -151.232, -151.2247, -151.1937, -151.1926, -151.1784, -151.1785, 
    -151.1404, -151.1555, -151.1236, -151.1622, -151.1496, -151.1489, 
    -151.1676, -151.2811, -151.3745, -151.4464, -151.4214, -151.4008, 
    -151.4007, -151.4126, -151.4712, -151.4349, -151.4413, -151.4486, 
    -151.4121, -151.4113, -151.444, -151.4505, -151.4251, -151.4113, 
    -151.4407, -151.3973, -151.397, -151.4028, -151.3982, -151.3973, 
    -151.3914, -151.396, -151.398, -151.4175, -151.3959, -151.3878, 
    -151.4011, -151.3826, -151.3811, -151.3866, -151.3923, -151.3905, 
    -151.3929, -151.3772, -151.3665, -151.3814, -151.3139, -151.2399, 
    -151.2403, -151.1985, -151.1742, -151.1026, -150.9694, -150.9747, 
    -150.9752, -150.9673, -150.9835, -150.9878, -150.9883, -150.9836, 
    -150.9971, -151.0244, -151.0126, -151.0047, -151.033, -151.0131, 
    -151.0613, -151.0434, -151.0566, -151.0353, -151.0142, -151.0128, 
    -151.0128, -151.0758, -151.2729, -151.3945, -151.1858, -151.4388, 
    -151.4537, -151.4695, -151.4878, -151.2489, -151.4948, -151.4949, 
    -151.5352, -151.566, -151.5519, -151.5524, -151.5441, -151.5395, 
    -151.5423, -151.5265, -151.5321, -151.583, -151.5251, -151.544, 
    -151.5457, -151.6007, -151.6711, -151.5275, -151.6807, -151.6799, 
    -151.7588, -151.7504, -151.5801, -151.58, -151.5717, -151.5077, 
    -151.5291, -151.5288, -151.4734, -151.4718, -151.4704, -151.4895, 
    -151.4801, -151.4954, -151.4872, -151.4852, -151.4155, -151.4466, 
    -151.4024, -151.3891, -151.3101, -151.3108, -151.3106, -151.3104, 
    -151.3064, -151.3096, -151.3047, -151.3117, -151.3048, -151.3164, 
    -151.302, -151.3178, -151.3411, -151.3718, -151.3826, -151.3421, 
    -151.3424, -151.1824, -151.2547, -151.2455, -151.255, -151.2489, 
    -151.2501, -151.2433, -151.2439, -151.2473, -151.2322, -151.2522, 
    -151.2516, -151.2508, -151.2489, -151.2322, -151.249, -151.2479, 
    -151.2543, -151.2458, -151.2531, -151.25, -151.2575, -151.2472, 
    -151.2359, -151.248, -151.2385, -151.2384, -151.2564, -151.2562, 
    -151.2507, -151.2577, -151.2391, -151.2594, -151.2665, -151.2656, 
    -151.2581, -151.2569, -151.2557, -151.2564, -151.2556, -151.3225, 
    -151.2646, -151.2769, -151.2664, -151.2745, -151.276, -151.2752, 
    -151.2823, -151.2891, -151.2888, -151.2679, -151.2331, -151.2448, 
    -151.2831, -151.2517, -151.2539, -151.2538, -151.2546, -151.2497, 
    -151.2499, -151.2505, -151.2659, -151.2608, -151.2583, -151.2601, 
    -151.2486, -151.2595, -151.261, -151.2407, -151.2428, -151.238, 
    -151.2563, -151.3509, -151.3448, -151.34, -151.2362, -151.3222, -151.328, 
    -151.3396, -151.3333, -151.3503, -151.379, -151.3628, -151.3611, 
    -151.353, -151.3678, -151.3404, -151.3401, -151.3602, -151.3577, 
    -151.3559, -151.361, -151.3966, -151.3951, -151.3587, -151.3591, 
    -151.3594, -151.3635, -151.3613, -151.3593, -151.3607, -151.361, 
    -151.3481, -151.3851, -151.415, -151.4486, -151.4363, -151.4312, 
    -151.4746, -151.4573, -151.4735, -151.4952, -151.4749, -151.4762, 
    -151.5246, -151.5407, -151.4763, -151.4767, -151.5583, -151.5625, 
    -151.5904, -151.5653, -151.608, -151.641, -151.5674, -151.6527, 
    -151.6458, -151.6573, -151.6544, -151.6599, -151.6578, -151.66, -151.664, 
    -151.6496, -151.6645, -151.6655, -151.6658, -151.6376, -151.7105, 
    -151.6395, -151.6829, -151.6351, -151.605, -151.5947, -151.5724, 
    -151.5694, -151.4315, -151.4175, -151.5792, -151.406, -151.3878, 
    -151.4032, -151.3738, -151.3718, -151.3555, -151.3626, -151.3593, 
    -151.3188, -151.364, -151.3598, -151.3602, -151.3335, -151.3714, 
    -151.3561, -151.36, -151.3922, -151.3592, -151.3598, -151.3733, 
    -151.3188, -151.3385, -151.3575, -151.3612, -151.3594, -151.3527, 
    -151.3485, -151.3833, -151.1943, -151.2452, -151.2523, -151.2353, 
    -151.2482, -151.251, -151.2448, -151.2538, -151.2678, -151.247, 
    -151.2545, -151.2472, -151.2484, -151.2477, -151.2479, -151.242, 
    -151.2375, -151.2474, -151.1986, -151.1282, -151.1287, -151.1761, 
    -151.1405, -151.1392, -151.1661, -151.1702, -151.1683, -151.1202, 
    -151.0326, -151.0189, -151.0282, -150.9467, -151.0338, -150.9965, 
    -150.9485, -150.9871, -150.9807, -150.9896, -150.9985, -150.9932, 
    -151.0177, -150.9987, -150.9993, -151.0199, -151.0279, -151.0337, 
    -150.9797, -151.0155, -151.0163, -151.0166, -151.0027, -151.014, 
    -151.0231, -151.0168, -151.0288, -151.0308, -150.9787, -150.9777, 
    -151.0402, -150.9674, -150.9401, -150.9946, -151.0221, -150.9881, 
    -151.0355, -151.0088, -151.0309, -151.0091, -150.9758, -151.048, 
    -150.9855, -150.9989, -151.033, -151.0019, -151.0146, -151.0186, 
    -151.0197, -151.0152, -151.0195, -151.0334, -151.0236, -151.0312, 
    -151.0254, -150.9946, -151.0269, -151.0282, -150.9949, -151.1, -151.1507, 
    -151.1554, -151.1964, -151.2004, -151.2826, -151.32, -151.299, -151.2935, 
    -151.2745, -151.2715, -151.3105, -151.3189, -151.3206, -151.3288, 
    -151.3351, -151.3067, -151.3649, -151.3411, -151.3531, -151.3038, 
    -151.3037, -151.3037, -151.2819, -151.2283, -151.2235, -151.1026, 
    -151.1526, -151.081, -151.2104, -151.021, -151.0175, -151.2051, 
    -151.0208, -151.031, -151.1419, -151.147, -151.1358, -151.0457, 
    -150.9921, -151.0306, -151.0266, -150.9916, -150.9912, -150.9752, 
    -150.9759, -150.9633, -150.9437, -150.9495, -150.963, -151.0283, 
    -151.0323, -150.9897, -150.9709, -150.9007, -150.9706, -150.9745, 
    -150.9868, -150.9916, -151.0063, -151.0047, -151.0185, -151.022, 
    -151.027, -151.0263, -151.0171, -151.0163, -151.0229, -151.1281, 
    -151.0446, -151.0365, -151.3953, -151.3987, -151.436, -151.4169, 
    -151.5211, -151.5202, -151.47, -151.5632, -151.3622, -151.362, -151.6454, 
    -151.3555, -151.3252, -151.5031, -151.5059, -151.5033, -151.5031, 
    -151.5188, -151.5074, -151.5316, -151.5379, -151.4891, -151.5472, 
    -151.5715, -151.5521, -151.5569, -151.5657, -151.5608, -151.5623, 
    -151.5937, -151.5784, -151.5667, -151.4439, -151.4323, -151.414, 
    -151.3832, -151.7393, -151.4206, -151.4505, -151.6701, -151.7018, 
    -151.5618, -151.5668, -151.5971, -151.5667, -151.5582, -151.5753, 
    -151.5955, -151.6116, -151.6307, -151.6428, -151.5987, -151.5697, 
    -151.6382, -151.6325, -151.6255, -151.6586, -151.6644, -151.6623, 
    -151.6509, -151.6587, -151.6599, -151.6565, -151.6597, -151.6572, 
    -151.6558, -151.6558, -151.6585, -151.6513, -151.6651, -151.6673, 
    -151.6555, -151.6596, -151.6587, -151.6628, -151.6524, -151.6596, 
    -151.6625, -151.6704, -151.6621, -151.6532, -151.6648, -151.6435, 
    -151.4607, -151.468, -151.4675, -151.466, -151.4737, -151.4585, -151.467, 
    -151.4867, -151.4762, -151.4753, -151.4707, -151.4683, -151.4698, 
    -151.4746, -151.4756, -151.4838, -151.5059, -151.5243, -151.4702, 
    -151.4666, -151.461, -151.4523, -151.4464, -151.4391, -151.3701, 
    -151.3575, -151.3636, -151.361, -151.3476, -151.3452, -151.3491, 
    -151.3316, -151.3281, -151.3249, -151.3287, -151.3549, -151.3649, 
    -151.3786, -151.3705, -151.3647, -151.3681, -151.3719, -151.3699, 
    -151.3664, -151.3635, -151.3575, -151.3573, -151.3505, -151.3625, 
    -151.2993, -151.3671, -151.3688, -151.3694, -151.2719, -151.3665, 
    -151.3613, -151.362, -151.3614, -151.3394, -151.3426, -151.3513, 
    -151.3564, -151.3439, -151.3973, -151.408, -151.3675, -151.3542, 
    -151.3572, -151.1804, -151.1823, -151.3062, -151.3729, -151.439, 
    -151.3317, -151.3397, -151.3379, -151.3284, -151.3378, -151.3294, 
    -151.3481, -151.3301, -151.3363, -151.3254, -151.3369, -151.3361, 
    -151.3367, -151.3356, -151.3366, -151.3465, -151.3443, -151.3575, 
    -151.354, -151.3516, -151.3565, -151.3669, -151.3663, -151.3893, 
    -151.3714, -151.3875, -151.4362, -151.4633, -151.4518, -151.3585, 
    -151.2643, -151.2583, -151.277, -151.3963, -151.2989, -151.2989, 
    -151.3195, -151.3329, -151.3221, -151.2772, -151.2812, -151.2979, 
    -151.2751, -151.2919, -151.255, -151.2894, -151.2636, -151.2412, 
    -151.2298, -151.218, -151.2404, -151.243, -151.2408, -151.2419, 
    -151.2419, -151.2365, -151.2388, -151.3542, -151.3846, -151.2494, 
    -151.4814, -151.5053, -151.6018, -151.6021, -151.6184, -151.626, 
    -151.6358, -151.6448, -151.6493, -151.6647, -151.6601, -151.6583, 
    -151.6622, -151.6591, -151.6618, -151.6661, -151.6635, -151.6629, 
    -151.6572, -151.6598, -151.6518, -151.6614, -151.6628, -151.6706, 
    -151.676, -151.6631, -151.66, -151.6543, -151.6587, -151.6628, -151.6349, 
    -151.7274, -151.5672, -151.5715, -151.5966, -151.5608, -151.5684, 
    -151.5546, -151.5474, -151.5366, -151.4895, -151.5155, -151.5042, 
    -151.4758, -151.4685, -151.4583, -151.4471, -151.4945, -151.4457, 
    -151.4574, -151.4883, -151.4398, -151.4041, -151.3469, -151.3101, 
    -151.2922, -151.3051, -151.2675, -151.267, -151.2626, -151.2714, 
    -151.2635, -151.2385, -151.2403, -151.2032, -151.1895, -151.2402, 
    -151.2366, -151.2373, -151.2444, -151.2469, -151.2473, -151.2508, 
    -151.2297, -151.1831, -151.2234, -151.2476, -151.2461, -151.2416, 
    -151.2283, -151.2419, -151.2376, -151.2802, -151.2543, -151.2487, 
    -151.1952, -151.2808, -151.2963, -151.3214, -151.3332, -151.1847, 
    -151.1904, -151.3755, -151.1764, -151.1921, -151.3107, -151.2923, 
    -151.2917, -151.3069, -151.3026, -151.306, -151.3006, -151.2195, 
    -151.2182, -151.2448, -151.2473, -151.2416, -151.2178, -151.2217, 
    -151.0991, -151.0793, -151.2456, -151.1799, -151.0374, -151.0546, 
    -151.0521, -151.241, -151.3364, -151.3813, -151.362, -151.3565, 
    -151.3639, -151.3522, -151.3587, -151.3643, -151.4011, -151.4021, 
    -151.4211, -151.3673, -151.4132, -151.419, -151.4684, -151.4148, 
    -151.4178, -151.4171, -151.4186, -151.4309, -151.4305, -151.4319, 
    -151.4331, -151.4351, -151.4454, -151.4251, -151.4238, -151.4373, 
    -151.4548, -151.4511, -151.4523, -151.4519, -151.4389, -151.4495, 
    -151.4531, -151.4649, -151.4918, -151.5133, -151.4881, -151.4845, 
    -151.5626, -151.5504, -151.533, -151.5127, -151.5086, -151.4855, 
    -151.4242, -151.4156, -151.4315, -151.4285, -151.4228, -151.4244, 
    -151.4175, -151.4226, -151.4271, -151.4486, -151.4478, -151.4494, 
    -151.3985, -151.3881, -151.3862, -151.3825, -151.3823, -151.3543, 
    -151.3328, -151.3302, -151.3436, -151.328, -151.36, -151.3541, -151.3056, 
    -151.331, -151.309, -151.3141, -151.2747, -151.3084, -151.2224, 
    -151.2093, -151.2089, -151.1747, -151.188, -151.2061, -151.2555, 
    -151.1949, -151.193, -151.1876, -151.1882, -151.1895, -151.183, 
    -151.1932, -151.1886, -151.1972, -151.1882, -151.1896, -151.1877, 
    -151.1881, -151.1872, -151.1872, -151.1873, -151.1873, -151.1875, 
    -151.1942, -151.1878, -151.1838, -151.1874, -151.1926, -151.1921, 
    -151.1894, -151.19, -151.1863, -151.1781, -151.1749, -151.178, 159.0115, 
    -109.17, -151.2062, -151.2054, -151.2029, -154.258, -154.2539, -154.1962, 
    -151.1256, -153.9989, 160.9647, -151.052, -151.0473, -151.1043, 
    -151.0677, -151.1958, -151.2589, -151.2755, -151.2757, -151.2757, 
    -151.3457, -151.335, -151.3432, -151.361, -151.3805, -151.4404, -151.582, 
    -151.5995, -151.6461, -151.655, -151.636, -151.6605, -151.663, -151.6543, 
    -151.6512, -151.6565, -151.6552, -151.6751, -151.6615, -151.6623, 
    -151.6602, -151.6669, -151.6542, -151.6538, -151.6579, -151.6576, 
    -151.6727, -151.6654, -151.6578, -151.6553, -151.6539, -151.6569, 
    -151.6635, -151.6604, -151.6444, -151.6356, -151.6379, -151.6353, 
    -151.6416, -151.6463, -151.5834, -151.5986, -151.5791, -151.5783, 
    -151.5737, -151.4812, -151.5553, -151.436, -151.3451, -151.3355, 
    -151.4709, -151.335, -151.3359, -151.3655, -151.2626, -151.2642, 
    -151.3621, -151.3577, -151.3555, -151.3611, -151.3512, -151.3654, 
    -151.365, -151.3637, -151.3636, -151.3554, -151.3452, -151.3654, 
    -151.3652, -151.366, -151.3654, -151.3612, -151.3554, -151.3043, 
    -151.3042, -151.2965, -151.3027, -151.3049, -151.3069, -151.3001, 
    -151.3019, -151.3014, -151.3008, -151.2988, -151.3087, -151.3062, 
    -151.3067, -151.3112, -151.3032, -151.2902, -151.2937, -151.3091, 
    -151.3278, -151.3169, -151.3168, -151.3303, -151.3204, -151.3249, 
    -151.3135, -151.3192, -151.3099, -151.3295, -151.2998, -151.2904, 
    -151.3131, -151.3741, -151.4212, -151.4446, -151.4446, -151.4402, 
    -151.2924, -151.2287, -151.2294, -151.2293, -151.2495, -151.2487, 
    -151.2369, -151.2414, -151.2542, -151.2656, -151.2501, -151.2635, 
    -151.261, -151.228, -151.2421, -151.2433, -151.2402, -151.2472, 
    -151.2401, -151.2451, -151.2401, -151.2473, -151.2476, -151.2455, 
    -151.2535, -151.2694, -151.2563, -151.2202, -151.3241, -151.3221, 
    -151.3503, -151.3547, -151.3503, -151.4299, -151.4897, -151.4972, 
    -151.509, -151.5262, -151.5358, -151.5452, -151.5518, -151.3552, 
    -151.6626, -151.6792, -151.6656, -151.656, -151.648, -151.6616, 
    -151.6405, -151.6595, -151.6951, -151.6613, -151.6585, -151.661, 
    -151.6595, -151.6647, -151.6647, -151.6574, -151.6392, -151.645, 
    -151.6277, -151.6466, -151.7159, -151.6754, -151.6768, -151.6108, 
    -151.5586, -151.5523, -151.5508, -151.5137, -151.4156, -151.4992, 
    -151.4156, -151.3997, -151.4326, -151.4073, -151.4022, -151.3794, 
    -151.3789, -151.3814, -151.3591, -151.3577, -151.3078, -151.3105, 
    -151.3085, -151.3128, -151.3187, -151.3036, -151.3052, -151.2906, 
    -151.318, -151.2731, -151.3104, -151.3116, -151.3123, -151.3317, 
    -151.3386, -151.3418, -151.3253, -151.3175, -151.3131, -151.3485, 
    -151.346, -151.3401, -151.3412, -151.3484, -151.3415, -151.3459, 
    -151.3588, -151.2507, -151.351, -151.3508, -151.3544, -151.3573, 
    -151.334, -151.3576, -151.3652, -151.3332, -151.3383, -151.3549, 
    -151.3173, -151.3378, -151.3398, -151.32, -151.3925, -151.4655, 
    -151.6608, -151.4035, -151.4253, -151.4014, -151.4064, -151.3985, 
    -151.4282, -151.4274, -151.4267, -151.4271, -151.4269, -151.4756, 
    -151.4755, -151.484, -151.5298, -151.504, -151.518, -151.5293, -151.5341, 
    -151.5555, -151.573, -151.5728, -151.6729, -151.5309, -151.421, 
    -151.4201, -151.4182, -151.4259, -151.4202, -151.4335, -151.4344, 
    -151.4167, -151.4131, -151.3442, -151.3339, -151.4201, -151.4182, 
    -151.3983, -151.3209, -151.3186, -151.32, -151.4089, -151.4002, 
    -151.4007, -151.3904, -151.4385, -151.4017, -151.4675, -151.4798, 
    -151.5172, -151.4962, -151.5376, -151.5589, -151.5496, -151.5576, 
    -151.5415, -151.6378, -151.6263, -151.6465, -151.6203, -151.536, 
    -151.3406, -151.4375, -151.7052, -151.4933, -151.4689, -151.4549, 
    -151.4543, -151.4326, -151.4528, -151.4584, -151.4446, -151.5005, 
    -151.4902, -151.5011, -151.5066, -151.5092, -151.513, -151.5176, 
    -151.4979, -151.5344, -151.5179, -151.5499, -151.5166, -151.5204, 
    -151.5145, -151.5203, -151.6127, -151.6711, -151.7838, -151.7567, 
    -151.6602, -151.6593, -151.6516, -151.6555, -151.6554, -151.6564, 
    -151.6564, -151.6446, -151.6277, -151.6307, -151.5713, -151.5624, 
    -151.5634, -151.5641, -151.5292, -151.5591, -151.5556, -151.5083, 
    -151.4928, -151.4859, -151.5441, -151.5403, -151.5336, -151.5347, 
    -151.5351, -151.4585, -151.5079, -151.4827, -151.4754, -151.4785, 
    -151.4327, -151.433, -151.4301, -151.4276, -151.4268, -151.4292, 
    -151.423, -151.4037, -151.404, -151.4305, -151.4306, -151.3848, 
    -151.4453, -151.3586, -151.435, -151.4391, -151.472, -151.4659, 
    -151.4627, -151.4534, -151.4611, -151.4598, -151.4488, -151.4492, 
    -151.3666, -151.3511, -151.3638, -151.3391, -151.3259, -151.3382, 
    -151.3223, -151.3352, -151.3257, -151.3197, -151.282, -151.2725, 
    -151.2533, -151.2641, -151.2687, -151.2555, -151.235, -151.2298, 
    -151.2353, -151.238, -151.2419, -151.2086, -151.2085, -151.1931, 
    -151.1755, -151.1764, -151.1931, -151.1938, -151.1933, -151.1896, 
    -151.1902, -151.1809, -151.1991, -151.1856, -151.181, -151.1872, 
    -151.1904, -151.1904, -151.2196, -151.2196, -151.2077, -151.2331, 
    -151.2094, -151.2603, -151.2733, -151.242, -151.2053, -151.1974, 
    -151.2086, -151.2298, -151.3522, -151.4041, -151.4031, -151.3785, 
    -151.4048, -151.4214, -151.4356, -151.4289, -151.429, -151.4269, 
    -151.4252, -151.6214, -151.4807, -151.4274, -151.4272, -151.481, 
    -151.4305, -151.4425, -151.4274, -151.4316, -151.4473, -151.4429, 
    -151.4403, -151.4312, -151.4407, -151.4361, -151.4378, -151.4593, 
    -151.4488, -151.4457, -151.4511, -151.4548, -151.4482, -151.4497, 
    -151.4317, -151.4503, -151.4535, -151.4587, -151.4572, -151.4971, 
    -151.4485, -151.4733, -151.4763, -151.6194, -151.685, -151.6637, 
    -151.6566, -151.6598, -151.6665, -151.671, -151.6427, -151.6405, 
    -151.6401, -151.6289, -151.6082, -151.63, -151.5935, -151.6247, 
    -151.6183, -151.6184, -151.5379, -151.5993, -151.5979, -151.5941, 
    -151.3882, -151.3931, -151.3273, -151.3135, -151.289, -151.2858, 
    -151.2673, -151.2592, -151.2534, -151.2414, -151.2443, -151.2455, 
    -151.2463, -151.248, -151.2473, -151.2443, -151.2446, -151.245, -151.244, 
    -151.2303, -151.2274, -151.2324, -151.2363, -151.2298, -151.2061, 
    -151.2409, -151.2447, -151.2307, -151.2306, -151.226, -151.2325, 
    -151.0817, -151.2759, -151.2775, -151.2444, -151.2711, -151.2371, 
    -151.2525, -151.1992, -151.199, -151.1808, -151.1721, -151.1615, 
    -150.9772, -151.3657, -151.3782, -151.4226, -151.4158, -151.4048, 
    -151.4465, -151.4547, -151.4733, -151.4157, -151.4212, -151.472, 
    -151.4484, -151.4233, -151.4215, -151.4312, -151.4329, -151.4417, 
    -151.4392, -151.4212, -151.4287, -151.4456, -151.4277, -151.4463, 
    -151.4443, -151.4456, -151.483, -151.494, -151.5026, -151.4844, 
    -151.5526, -151.648, -151.6296, -151.6609, -151.6605, -151.6608, 
    -151.6626, -151.6531, -151.6637, -151.6571, -151.6571, -151.6468, 
    -151.7162, -151.6091, -151.6154, -151.6193, -151.456, -151.5848, 
    -151.4286, -151.4298, -151.4292, -151.4299, -151.4299, -151.4295, 
    -151.4271, -151.4296, -151.4065, -151.4297, -151.4266, -151.4266, 
    -151.4162, -151.414, -151.4179, -151.4152, -151.4129, -151.4462, 
    -151.4455, -151.4333, -151.429, -151.4289, -151.3976, -151.4335, 
    -151.4291, -151.4221, -151.4191, -151.4226, -151.3955, -151.4083, 
    -151.4132, -151.3863, -151.4114, -151.4184, -151.4299, -151.4303, 
    -151.4301, -151.3977, -151.379, -151.3629, -151.3028, -151.3053, 
    -151.2835, -151.2756, -151.2757, -151.2688, -151.2707, -151.1789, 
    -151.1864, -151.1875, -151.1867, -151.2176, -151.2429, -151.2503, 
    -151.2583, -151.2383, -151.4204, -151.4244, -151.5096, -151.5277, 
    -151.5489, -151.2589, -151.5228, -151.5449, -151.5535, -151.5546, 
    -151.5388, -151.5552, -151.5323, -151.5357, -151.5314, -151.5395, 
    -151.5475, -151.5935, -151.6052, -151.6129, -151.6216, -151.6415, 
    -151.63, -151.6552, -151.6596, -151.7233, -151.6477, -151.6603, 
    -151.6524, -151.6723, -151.6593, -151.6616, -151.7825, -151.6833, 
    -151.6789, -151.6316, -151.632, -151.6364, -151.6339, -151.6386, 
    -151.6366, -151.6601, -151.6641, -151.664, -151.6544, -151.6374, 
    -151.625, -151.6138, -151.6041, -151.5863, -151.6365, -151.6178, 
    -151.5733, -151.5645, -151.556, -151.551, -151.5668, -151.5618, 
    -151.5653, -151.5675, -151.5356, -151.566, -151.5632, -151.4328, 
    -151.5402, -151.4146, -151.4147, -151.4313, -151.3954, -151.4716, 
    -151.3913, -151.4208, -151.4088, -151.4102, -151.4131, -151.4219, 
    -151.4386, -151.4482, -151.4485, -151.4489, -151.4486, -151.4837, 
    -151.4906, -151.487, -151.4954, -151.5233, -151.5593, -151.6049, 
    -151.5893, -151.6222, -151.6415, -151.6614, -151.6629, -151.7345, 
    -151.6374, -151.6957, -151.6528, -151.66, -151.6655, -151.6314, 
    -151.5942, -151.653, -151.6528, -151.6638, -151.6613, -151.619, 
    -151.6457, -151.5944, -151.6311, -151.5466, -151.5017, -151.4646, 
    -151.4474, -151.4296, -151.429, -151.4343, -151.4283, -151.4304, 
    -151.4296, -151.425, -151.4082, -151.4306, -151.4246, -151.4253, 
    -151.433, -151.4225, -151.4242, -151.4335, -151.4171, -151.4148, 
    -151.4043, -151.4309, -151.4281, -151.425, -151.4247, -151.4261, -151.42, 
    -151.4482, -151.5269, -151.5176, -151.5182, -151.5223, -151.5208, 
    -151.5235, -151.6574, -151.6587, -151.6641, -151.6739, -151.6516, 
    -151.6595, -151.6674, -151.6634, -151.6673, -151.6661, -151.6667, 
    -151.6518, -151.6608, -151.6606, -151.6593, -151.6597, -151.6579, 
    -151.6648, -151.6577, -151.6634, -151.6365, -151.5863, -151.65, 
    -151.6499, -151.6588, -151.6258 ;

 offset = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _ ;

 offset_orientation = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 platform = _ ;

 qartod_location_flag = _ ;

 qartod_rollup_flag2 = _ ;

 qartod_speed_flag = _ ;

 qartod_time_flag = _ ;

 semi_major_axis = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, 1729, 449, 1879, 4155, 896, 7131, 215, 698, 4728, _, _, _, _, _, _, _, 
    3950, _, _, 3629, _, 7713, _, _, 50071, 19560, 6071, 13584, _, 2509, 
    2749, _, 3542, _, 3830, 2202, 2684, _, _, 2654, _, _, 2953, _, _, 4394, 
    _, 5287, 7608, 5741, 6199, 2802, 2808, 29680, 4270, 3691, _, _, _, 7550, 
    _, 4711, _, 6220, 7789, 6262, 6292, 23300, 3373, 1317, 6878, 3268, 12331, 
    87186, 13782, 2710, 22882, 12692, 4208, 3938, 3939, 4081, 1574, 2901, 
    959, 2076, 2230, 4322, 3101, 2964, 5800, 1428, 1436, 33933, _, 4553, 
    4805, 8034, 1762, 4042, 4264, 8304, 58044, 5173, 1572, _, 1188, 1353, 
    748, 721, 2106, _, _, _, _, _, _, _, _, _, _, _, 646, 1222, 4598, 3061, 
    _, 3824, 598, 409, 2797, 30451, 7421, _, 6620, 7438, 5195, 2716, 2186, 
    438, 294, 563, 8033, 1425, 465, 1871, 590, 2047, 11150, _, _, _, _, _, _, 
    _, _, _, _, 483, _, _, _, 2147, 46278, 5551, 5044, 4681, 4722, 4452, 447, 
    34721, 11316, 3742, 2067, 6818, 4349, 3129, 2419, 1336, _, _, 2811, _, _, 
    _, 5212, 6213, 1798, 1915, 877, 2023, 3894, 1947, 1934, 1275, 743, 4553, 
    183, 2263, 571, 895, _, 1317, 2615, 3117, 29216, 45595, 147837, 39977, 
    14474, _, _, _, _, _, _, _, _, _, _, 8031, 1031, 1335, _, _, 31990, _, 
    4760, 2324, 991, 386, _, 784, 578, _, 1309, _, 1810, _, 808, 2459, 3272, 
    887, 1813, 31007, 1037, 479, 1611, 2976, 1493, _, _, 5514, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 15433, _, 100164, 14557, 
    14274, 9836, 1317, _, 2500, 1995, 13284, 7079, 4218, 717, 1711, 1465, 
    1766, 25816, 11744, 281, 2537, _, 7394, 5284, _, _, _, _, _, _, _, _, _, 
    _, 706, 1021, 519, 2265, 422, 386, 1775, 11668, 1334, 1679, 330, 1128, 
    526, 412, 676, 1985, 2111, 1532, 3089, 775, 1034, 1496, 1411, 2795, 
    70736, 103176, 708, 470, 2328, 2513, 2669, 12538, 12819, 5509, 728, 673, 
    _, 18456, _, _, 11311, 1344, 2457, _, 1161, _, 14575, 1584, 569, 3526, 
    1690, 1302, _, 5388, _, 13838, _, 5070, _, 3528, 2645, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, 4792, 54875, _, _, _, 13447, 2999, _, _, _, 
    _, 2182, _, 6981, 1783, _, 1047, 799, _, 1173, 455, _, 1480, 1588, 1794, 
    1933, 8479, 3550, _, 168109, 16987, 25699, _, 19019, 10778, 14590, _, _, 
    _, _, _, _, _, 71971, _, 5943, _, 1924, 31386, 409, 1179, 9862, 2303, 
    2259, 2451, 16082, 1751, _, _, _, _, 21987, _, _, 1341, _, 3053, _, 6593, 
    _, 7430, 2336, 2371, 6682, 15352, 4092, _, 7392, 3087, 5181, 2028, 14985, 
    3065, 2105, 948, 435, 2950, _, _, 3309, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, 1041, 4263, _, 21318, _, 4748, _, 
    13988, 1899, _, 3611, 2413, 15003, 4092, 1460, 1879, 389, _, _, _, 6409, 
    2018, _, _, 7989, _, 901, _, 674, 1074, 6349, 7392, _, _, _, _, _, _, _, 
    _, _, _, _, _, 103628, 36405, 4758, 1578, _, 1556, 20791, _, 2820, 2115, 
    620, 27583, 2904, 2530, 32131, 7651, 611, _, _, 2582, 13979, 1209, 1823, 
    540, 350, 16340, 163291, 37454, _, 649, 1252, 2023, 964, 4136, 52568, 
    26566, 4734, 41719, 11640, 899, 964, 705, 7878, 7916, 8325, 8194, _, _, 
    _, 55076, 9782, _, 249251, 28150, 15123, 12594, 2826, 1212, 1329, _, 
    2200, 305, 52663, 4189, 2566, 3151, 31595, 1486, 9548, 1401, 5031, _, 
    5299, 5062, 2309, _, _, _, _, _, _, _, _, 4572, _, _, _, _, _, 3396, _, 
    _, _, 9001, _, 3642, 2490, _, _, _, 3504, 49573, 13231, 1073, _, 9850, 
    2063, _, 2959, 8419, _, 9794, _, 11224, 711, _, _, _, _, 4727, 5898, _, 
    11785, _, 6448, _, _, _, _, 1050, _, 2793, _, _, _, _, 6550, 7698, 513, 
    6250, 943, 404, 562, 1952, 637, 288, 891, 2211, 2571, 4670, 2374, 1487, 
    505, 15653, 1121, 3660, 555, 2118, 4121, 1458, _, _, _, _, _, _, _, _, _, 
    _, 4331, 47509, 13052, _, _, 3157, _, 6697, 1280, 501, 5959, 615, 730, 
    39232, 1974, 467, 426, 2534, 578, 3128, 1084, 416, 529, 2284, 3556, _, _, 
    _, _, _, _, _, 23439, 16782, 15614, 193597, 1253, 2229, 1953, 1807, 568, 
    9193, 8591, 408, 715, 4074, 3330, _, 890, 1656, _, _, _, _, 6642, 4118, 
    _, 3339, _, 21094, 7492, 1367, 23198, 2332, 2007, 821, 1496, 854, 296, 
    826, 2588, 793, 570, 6402, 39285, 2598, _, _, 2838, _, _, 16189, 35592, 
    1586, 1017, 555, 336, 1392, 5749, 2144, 2257, 9051, 26000, 2250, 2457, 
    1749, 6370, 2276, 29303, _, _, _, _, 7091, 12715, 17308, 2549, 2461, 
    2785, 3058, _, _, 22951, 5895, 5927, _, 5500, _, _, 18725, 2009, 3773, 
    9177, _, 4152, 11904, _, 4398, 4771, _, 395, 1557, 1440, 503, 35664, 
    9450, 5256, 3163, _, _, 7591, 447, 557, 1627, 2134, 3707, _, 1294, 1335, 
    790, 2389, 582, 2832, 3520, 29232, 872, 1658, 3167, 6184, 1766, 2183, _, 
    _, 2874, _, _, _, _, _, _, _, 6340, _, 1652, 2354, 3209, _, 759, 1410, 
    4462, 4175, 1940, 497, 545, _, 5913, 8588, 2099, 1311, 1513, 2767, 649, 
    1827, 4725, 20261, 8403, 7910, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    714, 20096, 2574, 648, 3921, 2401, 561, 743, 3459, 455, 15741, 234, 473, 
    740, 4554, 1083, 2828, 4243, 7058, 2801, 13731, 29772, 222996, 12956, 
    10621, 11712, 10364, _, _, _, _, _, _, _, _, 6253, 2731, _, _, _, _, 
    1031, 303, 921, 918, 25053, 4564, 44344, 33106, 61765, 4714, 4876, 257, 
    1621, _, 2168, _, 3207, _, _, 4447, 32821, 3666, 3767, _, 3478, _, 1908, 
    1563, 2679, 5300, 7643, 1088, 57213, 3164, 42008, 2682, 73806, 1375, 
    4459, 471, 1368, 4766, _, 45254, 1545, _, _, 1706, 3755, 32595, 5071, 
    4689, 36937, 8981, 2980, 474, 220, 865, 212, 771, 2290, 1184, 1183, 1319, 
    1178, _, 2287, _, 184243, _, 3362, _, 450, _, 790, 1355, _, _, _, _, _, 
    11930, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, 567, _, 4036, _, _, 855, 1367, 1726, _, _, 1209, 1736, 459, 
    1051, _, 973, 513, _, _, 6751, 557, _, _, 877, _, 2021, _, 1968, 608, _, 
    6738, _, 2543, _, 1375, _, 3849, _, 2177, 1735, 4395, 9695, 15092, _, _, 
    _, _, _, _, _, 6325, 8340, 8097, 48207, 1681, 9407, 4600, 794, 4833, 337, 
    999, 22402, _, 5716, 1303, 6953, 55570, 1116, 285, 1292, 2110, _, 5195, 
    _, 1987, 1781, 2288, 2526, 5890, _, _, 7079, _, _, 6811, 6864, 16131, 
    18863, 30033, _, 34714, 5979, _, 17820, 14670, _, 68539, _, 14633, _, _, 
    _, _, 4096, _, _, _, _, 585, 9533, 3556, 5600, 21873, 526, 5151, 614, 
    1813, 1001, 541, 1866, 7344, 37212, 378, _, 1744, _, _, 2528, _, 6012, _, 
    _, _, _, _, 9606, 6889, 2512, _, _, _, _, _, _, 28788, 11244, 11320, _, 
    3456, _, 2046, _, _, _, 365, 420, 934, 998, 590, 1451, 1824, 995, 572, 
    941, _, 9141, 2202, 11127, 421, 368, 2262, _, _, 5628, _, _, _, 87398, _, 
    _, 9454, 1155, 584, 1055, 1939, 3875, 3040, 468, 2940, 7878, 618, 553, 
    1186, 8205, 5820, 952, 358, 4150, 11238, 3762, 7775, 16840, 70477, _, 
    20246, 5756, _, 4461, 2315, 1641, 947, 2029, _, 11614, _, _, 5729, 5327, 
    4922, 4408, _, _, _, _, _, 6620, 628, _, _, _, _, 35409, _, _, 13437, _, 
    _, _, 1278, 2493, _, 22832, _, 3458, 16046, 5177, 4469, 22703, 2928, 
    6714, _, 2113, 1917, _, _, 21006, _, 7722, _, 2491, _, _, _, _, _, 3309, 
    _, 24759, _, _, 3420, 2245, _, _, 1062, 873, 1016, 3019, 332, 751, 927, 
    1777, 1550, 7610, 4487, 10311, 6695, 6601, 9856, 3197, 2456, 1375, 306, 
    1465, 14048, _, 6836, 7487, 7205, 12901, 7259, 7989, 6757, 15913, 61103, 
    16367, 8662, 6436, _, 4750, 1524, 5796, 2696, 2085, 2537, 2416, 2842, 
    15942, 1885, _, 29471, 37508, 30009, _, _, _, 17033, 4215, _, 455, 734, 
    1772, 2910, 662, 8083, 3767, 1361, 14433, _, _, 154016, 2405, _, 6051, 
    7111, 3083, _, _, 3903, 5163, 3103, _, 20135, 305766, 22337, _, 9969, _, 
    4545, 6563, 4525, 2598, 987, 1458, 42972, 8314, 107494, 2969, 1163, 3146, 
    _, 11833, 5175, 2659, 7460, 912, 1017, 13018, 1188, 5697, 950, 1818, 
    23414, 6689, 426, 1320, 878, 3471, 2097, _, _, _, _, _, _, 21955, _, _, 
    _, _, 128249, 205835, 3997, 7456, 15598, 36373, 11186, _, _, 18174, 398, 
    19221, 1790, 1042, 1700, 1049, 1722, 4141, 5643, _, _, _, 2795, _, _, _, 
    _, _, _, _, _, _, _, _, _, 3342, 1961, _, 6748, 964, 1027, 779, 802, 
    2149, 6377, 14874, 1078, 1224, 1460, 1184, 647, 894, 2909, 15219, 273, 
    2436, _, _, 4257, 4836, 5957, 5924, 23428, 226506, 3110, 4570, 23908, 
    55857, 18969, 2233, 985, 4872, 1825, 1405, 4129, 3388, _, _, _, _, _, _, 
    6426, _, 1785, 6108, 8072, _, _, _, _, _, _, _, _, _, _, _, _, _, 5542, 
    514, 1352, 1527, _, 537, 18883, 2945, 5855, 8675, 2626, 18184, _, 6905, 
    1016, _, 1142, _, 1715, 11980, _, 6196, 561, _, _, 5422, 3775, _, 908, 
    1111, 2831, _, _, _, 10922, 14535, 13980, 12499, 1866, _, 15273, 2179, _, 
    2675, 2487, 2575, _, _, _, 241, 726, 2261, 13056, 2735, 1409, 1822, 677, 
    681, 3243, 448, 230, 3346, 457, 539, 474, 4176, 15179, 864, 1208, 1933, 
    656, 11656, _, 10368, _, _, _, _, 11867, _, _, 68196, _, 3764, 1537, 
    1819, 1942, 9916, 8298, 7851, 1429, _, 1372, 4779, 1788, 7690, 2148, 
    16404, _, _, 750, 2376, _, 12101, _, _, 10570, 7298, 3927, 1566, 1152, 
    2054, _, _, _, _, _, 11921, 2417, 3520, 3088, 254, 862, 13253, 557, 2158, 
    2647, 609, 3497, 2992, 666, 1080, 12938, 45201, _, 10691, 1097, 2361, 
    11545, 1761, 6324, 18564, _, _, _, _, _, _, _, _, _, _, 30383, 17230, 
    783, _, 1062, _, 2972, 1436, 13986, 8827, 912, 5475, 8841, _, 1044, 
    104255, 18250, 10469, 7109, 368, 15881, 3403, _, 499, 1761, 2195, 504, 
    11373, 4239, _, _, _, 16063, _, 8350, 11465, 4067, 125396, 2051, 2656, 
    3105, 3461, _, 18394, _, _, _, _, 7375, 9369, 9314, _, _, _, _, _, 1140, 
    1757, _, 4807, _, 295, 2531, 478, _, 880, 2144, 2044, 2060, 1623, 2288, 
    1463, 280, _, 1724, 3253, 1429, 5799, 1495, 4343, 8089, 4245, _, 268, 
    5469, 7869, _, 5732, 4218, 1552, 2043, 502, 303, 1114, 15174, 1387, 846, 
    454, 7904, 9450, 5546, 7188, 3124, 648, 1568, 3479, _, _, 13629, 443, 
    26104, 351, _, 1655, 1964, 1611, 1620, 38705, 637, 1413, 382, 2175, 439, 
    948, 1551, 30215, 4785, 416, 61904, 6856, 4775, 1123, _, _, _, 24518, _, 
    21008, 19971, 49090, 9220, _, 4373, 6849, 4755, 3446, _, _, 2454, 70492, 
    _, 2778, 85917, 7350, 8711, 6056, 3311, _, 4330, _, 40308, _, 897, _, 
    30229, 2342, 430, 3130, 3701, _, _, _, _, _, _, 7692, _, 18119, _, 12836, 
    843, _, _, 5780, _, 472, 1343, 581, 311, _, 3270, 2319, 53619, 2041, 
    2923, 454, _, 925, _, _, 1017, 1951, 3098, 1766, 28874, 10764, 3709, 
    2468, 1268, 13995, 10221, 1166, 647, _, _, _, _, _, _, _, _, _, _, _, 
    4220, 14399, _, 64595, 19295, _, 9353, 2905, 415, _, _, _, _, _, _, _, _, 
    _, _, 3249, _, _, 1851, _, 9860, 3438, _, 2451, _, 2609, _, 2916, 2926, 
    9003, _, 12809, _, 1655, _, 1591, _, _, 2355, 4317, 19840, 430, 822, 
    4997, 3889, 3466, _, 34726, _, _, 2014, 2309, 1214, 1745, 5801, _, 13918, 
    _, 622, 655, 1479, 338, 1161, 783, 4668, 2173, 176507, 2829, 504, 28344, 
    8605, 4371, 2225, 7421, _, _, 4536, 269, 990, 7491, 3709, 1471, 2187, 
    841, _, 2716, 3087, _, 377, 1531, 1139, 699, 1489, 1742, 3160, 1051, 
    8694, _, 52310, 1935, _, 1931, 2436, 2805, _, 4372, 519, _, _, _, _, 
    22155, _, 442, _, 1846, _, 8645, 13772, 557, 643, 1568, _, 8973, 4846, 
    27579, 1763, 1674, 2274, 26160, 2923, 499, 1692, 6399, 5529, 11885, 4555, 
    6709, _, _, _, _, _, 2266, _, 1860, 10752, 2909, 4553, _, _, _, _, _, _, 
    _, 5138, 3433, 3510, 394, 10880, 13776, 2670, 3744, _, 4653, 452, 2562, 
    273, 745, 3652, 101855, 3128, 4097, 1770, _, _, 1950, 2468, 1941, _, _, 
    _, _, _, 1104, 2923, 9351, 2322, _, 1669, 1824, 381, 7946, 953, 2260, 
    3561, 1030, 844, 1491, 1078, 540, _, _, 31232, 7305, 838, 14616, 13436, 
    3933, 1300, 1053, 1439, _, _, _, _, _, _, 435736, 16838, 18726, 997, 
    1589, 176029, 2449, 4940, 14093, 34902, 11613, 1580, 9837, 4640, _, 2438, 
    _, 2467, _, 647, _, _, _, _, _, _, _, _, 3040, 6562, 9265, 17347, _, _, 
    _, 11051, 16676, 73577, 65154, 25951, 53064, _, _, _, _, 186136, 4587, 
    2343, _, 18146, 14013, 6857, _, _, 682, 1845, 15388, 18010, _, 504, 355, 
    365, _, 13831, 3895, _, _, 8081, 39446, 4330, 3500, 1722, _, _, _, _, 
    3188, 3568, _, 16238, 2604, 1989, 2131, 2198, _, 3086, 3617, 3484, 6144, 
    1846, 2312, 22551, 3659, 5679, 1275, 1747, 1208, 432, 583, _, 679, 723, 
    _, _, _, 4403, _, _, _, 5579, _, 6762, _, 238, _, _, _, _, 7690, 4131, _, 
    1078, _, 3666, _, _, 28182, _, 16182, 1109, _, 1007, 1844, _, 2105, 2105, 
    2452, 3544, _, _, 26125, _, 5937, 6714, 8271, 6366, 472, 1051, 1542, 
    5891, 1489, 3426, 6172, 228666, _, 2835, _, 1462, 16937, 1856, _, _, 
    5807, 3685, _, 2116, 2253, _, _, _, 3177, 3381, 3545, 1544, 27631, _, _, 
    _, _, _, _, 4588, 9170, 279, 4852, 2911, 4073, 18637, 750, 1441, 5526, 
    6038, 1498, 1477, 3923, 3039, 41769, 1398, _, 37047, 998, 1168, 994, 
    1046, 493, 3467, 1795, _, _, _, 9911, 441, 3195, 300, 1088, 1557, 2062, 
    _, _, 258, 1065, 817, 520, 362, 6519, 999, 1679, 17204, 515, 13292, 6857, 
    2222, _, _, 13141, 554, _, 4279, 3613, _, 3456, 316, _, 3096, 4497, 1689, 
    22581, 1846, 3584, 3325, 3208, _, 6382, _, _, _, 7229, 7325, 26587, 
    11050, 7956, 1791, _, 2049, 1177, 1521, 2132, 5044, 1258, 511, _, 1719, 
    1949, 382, _, 3849, 2234, 1749, 386, _, 477, 4167, 3554, _, 273, 1551, 
    7134, 11104, _, _, _, _, 3649, 5114, _, _, _, 7656, _, _, 12777, 16141, 
    58905, 6903, _, _, _, 7308, _, _, 1973, _, 1821, 2170, _, 2742, _, _, 
    23626, _, _, 31867, 26391, _, 2268, 3474, _, 8624, 3222, _, 3943, 15894, 
    10326, 6454, 32437, _, 85617, _, 7773, 2013, _, 3631, 2264, 3543, 23491, 
    754, 863, 1560, 4685, 56509, 863, 894, _, 44911, 7637, _, 5280, 2935, 
    2575, _, 2218, _, 4494, _, _, _, _, _, _, _, 9869, 867, 45487, _, _, _, 
    _, 285, 2329, 3557, 5923, 134196, _, 5920, _, 19548, 727, 1193, 942, 
    1387, 1331, 4985, 881, 54970, 10553, 4043, 917, 1845, 972, 8844, 1221, 
    3828, _, _, _, _, _, _, _, 9791, 3492, 4348, 694, 5157, 23055, 720, _, 
    3193, 1111, _, _, 7794, 3986, 2769, _, 2253, 49357, 11522, 1026, 3008, _, 
    _, _, _, _, _, _, _, _, _, _, _, 27996, _, _, 27515, 4977, 5962, 7399, 
    3720, 5649, 4475, 3526, 3505, 609, 1795, 4043, 31698, 86199, 26736, 4938, 
    5705, 374, 925, 1358, 2324, 4373, 1474, 603, 284, 8115, 1219, 2345, 773, 
    532, 1392, 666, 759, 1163, 2861, 1857, 2191, 2108, 2744, 2821, 1090, 312, 
    2167, 3370, 4256, 616, 12035, 34094, _, _, _, _, _, _, _, _, _, _, 2418, 
    867, 487, 551, 1151, 3452, 1648, _, 4286, 1572, 3179, 5273, 23755, 402, 
    410, 1895, 2199, 1878, 359, 817, _, 351, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, 5322, 17964, _, _, 11807, _, _, 8632, 46985, 25442, 4124, 7198, 
    987, 434, 481, 25281, 471, 1847, 598, 5674, 2288, 1277, 715, 1580, 5130, 
    590, 9447, 8181, 610, _, 3081, 3515, _, _, _, _, _, _, 8889, _, 29943, _, 
    84009, 27626, 3270, 3724, _, 4370, 3842, _, 16121, 11786, _, 12786, _, 
    3289, _, 1483, _, 1854, 566207, 13862, _, 18363, 16881, 18592, 19046, 
    2930, 2938, _, _, _, _, _, 17338, _, _, 5391, 14133, _, _, 6194, 34266, 
    3152, 2141, 6715, 2786, 1863, 645, 1125, 1896, 1763, 1953, 12458, _, _, 
    _, _, _, _, _, 8585, 3363, _, _, 3628, 681, 2021, 937, 1367, 4752, _, 
    21210, 6354, 2126, 8824, 28770, _, 3702, _, 3454, _, _, 1121, 1214, _, 
    3760, 28850, _, _, _, _, 4796, 324, 749, 48130, 493, 994, 407, 439, 581, 
    647, 911, 991, 524, 643, 210, 1705, 1189, 6305, 383, 420, 4328, 4712, 
    8581, 345, 2438, _, _, _, 10154, _, 416, _, 2539, 7254, 3523, 4160, 7346, 
    107224, 4171, _, 5841, 779, 339, 1629, 1403, 5620, _, 44498, 27280, 4399, 
    1715, 3603, 4315, 2811, 2951, _, _, _, _, _, _, _, _, _, _, 44061, 973, 
    _, 632, 3289, 7115, 466, _, 5863, 4574, _, 6219, 12777, 7494, 2878, 5968, 
    756, 4256, 8808, _, 4126, 8202, _, 720, 932, _, _, _, _, _, _, _, _, _, 
    8598, 459, 6831, 7295, _, 6174, _, 1362, _, 3211, 2491, 1566, _, 13002, 
    2586, 2564, _, 213, 1400, 882, 6911, 5307, 4665, 8266, 6523, _, 34580, _, 
    868, 507, 1368, 1992, 13648, _, 17139, _, _, _, _, _, 23091, _, 43518, _, 
    _, _, _, _, _, _, _, _, 27548, 948, 582, 1918, 3774, 441, _, 401, _, _, 
    8130, 1374, 2855, 2246, _, _, 5805, 320, _, 1691, 17057, _, _, 1692, _, 
    3502, 2630, 13885, 3444, 1699, 2184, 2384, _, _, 37146, 4424, 2595, 7948, 
    5510, 1125, 4873, 1630, 1643, _, 3438, _, _, 3650, 11305, 2685, 814, 777, 
    1762, 5425, 1359, 1377, 1790, 573, 3773, 1431, 2013, 2606, _, 7456, _, 
    10775, 4436, _, _, _, 3363, 3994, 4369, 4630, 2578, 745, 4002, 2915, 
    3071, 1367, 3394, 3778, 3752, 3219, 7075, 9999, 5253, 34130, 6067, _, 
    4232, 4183, 1924, 1841, 3692, _, _, _, _, _, _, _, _, 59462, 42114, _, 
    26774, _, _, _, 140107, 16530, 6765, 6525, _, 4452, 3459, 8318, 369, 490, 
    1137, 266, 3063, 3783, 969, 12730, 2588, 3026, _, _, 3195, 3953, 3905, 
    371, _, 4690, 5397, _, _, 10926, 1776, 16205, 6974, 12150, 7355, 8106, 
    984, 5220, 1496, _, 5278, 1164, 311, 2416, 6449, 2631, 2014, 1208, 6753, 
    13600, 2508, 9917, 4440, 6525, 1160, 787, 285, _, _, _, _, _, _, 11824, 
    127873, 50086, _, _, 1973, 69706, _, _, 226543, 880, 671, 544, _, 4884, 
    _, _, 15958, _, 27883, 8947, _, 349, 7167, _, 4236, _, 1071, 3025, _, _, 
    _, _, _, _, _, _, _, 14492, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    7883, 92921, _, _, 11812, _, 6103, _, 1473, 802, 1947, 4118, 10341, 6850, 
    6903, 10399, 160751, 884, 2896, 9103, 30122, _, 21347, 2923, 1078, 1711, 
    1977, _, 4351, _, _, 714, _, 552, 1193, 1991, 849, 1599, 3405, 3701, 855, 
    15481, 9716, _, 9726, 1249, 506, 1924, _, _, 3755, 1657, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, 2891, _, _, 1568, 3210, 2844, 1425, 1921, 
    2278, 2076, 2535, 2817, 2947, 27223, 1379, 826, 597, 7113, 3684, 14054, 
    5065, _, 9936, _, _, _, _, 1218, 19038, 1072, 1810, 1944, 1908, 194, 
    1374, _, 1849, 6536, 641, 476, _, _, 467, 329, 7645, _, 291, _, _, 1835, 
    484, 1003, 1666, 411, 524, 5941, _, 1533, _, _, 5761, 441, _, _, 4639, _, 
    12262, 662, 856, 839, 609, 1071, 381, 297, 657, 2321, 257, 3162, 630, 
    1035, 10301, 5491, _, 1512, 3764, 7773, _, 9227, 7612, 619, 382, 1156, 
    2989, 3550, 2460, 2258, 35925, _, _, 4189, _, 4079, 4095, _, 4164, 19154, 
    2411, _, 1861, _, 1997, 2779, 3966, 581, 1081, 1225, 1789, 13937, 3917, 
    1407, 1696, 1266, 1186, 1900, 5498, 47289, 4047, 1208, 1667, 7489, 4701, 
    4354, 476, 661, 2041, 1506, 2456, _, _, 4820, 44252, 3471, 2015, 43883, 
    2912, _, _, _, 2706, 2806, 1165, 1528, 1568, 2114, 21703, 14321, 30306, 
    18822, 16186, 3443, 777, 2439, 1264, 1534, 628, _, 1036, 3974, 460, 254, 
    602, 21449, 7255, 4011, 2741, 2771, 2657, _, 19505, _, _, _, 7482, 83969, 
    34963, 13051, _, 1058, _, 33113, _, 3470, 1558, 2992, _, 5392, 1853, 
    8061, 2856, 66455, 52138, 31901, 4368, 1262, _, _, _, 5542, _, _, 176776, 
    _, _, _, _, 21188, 14986, 6292, 29038, _, 921, 1703, 327, 1236, 1764, _, 
    _, 1680, 481990, 12749, 15537, 7843, 566, 289577, 28731, _, 17348, 5027, 
    1358, 399, 585, 28995, 14167, 12986, 2059, 469, 436, 1660, 2509, 2875, 
    3905, 4861, 20035, 3400, 4011, 3583, _, _, _, _, 14149, 384, 1534, 3264, 
    649, 309, _, _, _, _, 4502, 15695, 15003, 1490, 1543, 3990, 5011, 5722, 
    310, 384, 405, _, 205357, 1458, 5562, 1522, 2792, 5035, 316, 5231, 6549, 
    _, 892, 3032, 767, _, 3942, _, 4512, 3357, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, 9373, _, _, _, 2704, _, 1491, _, 2081, 1506, _, 12276, 1705, 
    3807, 481, 2133, 4921, 13151, 507, 1990, 607, 1069, 550, 1604, 153, 9442, 
    533, 1742, 365, 1553, 1450, _, _, _, _, 20576, _, 785, _, 3583, 13454, 
    2037, 451, 1565, 273, 303, 12410, 4990, 388, 708, 974, 199, 72516, 
    129573, 825, 359, 1464, 1202, 351, 4342, _, _, _, _, _, _, _, _, 2980, _, 
    48498, _, 7823, 4913, _, _, 6650, 6877, 1150, _, _, 10470, 4566, _, 
    14900, _, 12324, 1716, 4897, _, 874, _, 1033, 831, 2349, 2765, 3519, _, 
    24234, _, 5421, _, _, 1253, 1946, 2254, _, _, 84066, _, _, 4325, 12269, 
    _, 9927, _, _, 8165, 282, _, _, 5405, 1062, 2848, _, 26676, _, _, 35104, 
    14693, 33753, 8333, 4374, _, _, _, 2091, 7179, _, 31814, 6275, _, 1275, 
    563, 638, 706, _, 2022, _, _, _, 4353, 8392, _, 2561, 3418, 21486, 14626, 
    _, 123239, 3118, _, _, _, 2922, 4527, _, _, 3890, _, _, 1065, _, 1279, _, 
    1640, _, 42307, 4208, 3753, 3795, 51851, 1987, 2179, 3475, 2109, 2003, 
    8666, 2153, _, _, _, _, 9811, 8978, _, 3764, 4523, 3522, _, 3784, _, 
    1608, _, 884, 54861, 4197, 71636, 60029, 23997, 576, 25226, 3905, 394, _, 
    1436, 2477, _, _, _, 16285, _, _, 2505, 2069, 4249, 1336, 1281, _, _, _, 
    _, _, _, 1417, _, 5762, 2963, 2237, _, _, 40848, 10809, 13759, 13321, 
    4010, 4076, 3054, 8644, 18833, _, 20468, _, 6041, _, _, 4699, _, _, 
    42986, 23321, 8880, 27141, _, 3700, 4369, 415, 712, 3423, 1542, _, 5720, 
    726, _, _, _, _, _, 4570, _, 18347, _, 972, 940, 497, 8701, 6493, 13713, 
    12040, 13781, 3006, 13967, _, 5533, 6750, _, 3905, 7610, 21147, 20824, 
    20468, 58379, 18039, 771, 2897, 27813, 1464, 1248, 1264, 993, 4261, 580, 
    1244, 27711, 9111, 4638, 1485, 616, 32580, _, 6809, 4818, 1110, 1002, 
    2025, 5780, 7461, _, _, _, _, 6773, _, _, 31048, 34920, 17998, 2308, 
    8382, 1326, 12126, 1981, _, _, _, _, 20425, 2251, _, 5918, 4083, 970, 
    258, 5030, 640, 487, 810, 371, 1383, 1153, 428, 428, 719, 949, 396, 397, 
    580, 10012, 337, 596, 14587, 3336, 4770, 1440, 676, 389, 9552, 8772, _, 
    1213, 1099, 3958, 72119, 592, _, 20714, 1283, 1376, 5021, 1871, 2095, 
    11966, 9819, 4343, 8289, 9518, 1224, 1328, 2066, 12350, _, 4235, 7710, _, 
    5148, 475, _, _, 26132, 20577, 3815, 5507, 1270, 966, 5168, 525, _, 1111, 
    3388, 4989, 34266, 3505, 19808, 359, 996, 2245, _, 8509, _, _, _, 13054, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, 23014, 110031, _, 157320, 
    25611, 1884, 1485, 810, 1947, 374, 1455, 1935, 1366, _, 910, 1670, _, _, 
    428, _, 3938, _, 1274, 3061, _, 5625, 41777, 2506, 3892, _, _, 6923, _, 
    31816, _, _, _, _, 4189, 5073, 4826, 1258, 1707, 1979, 4972, _, 1172, _, 
    2416, _, 1153, 2413, 603, 2577, 1692, _, 1067, 1200, 8568, 9605, 30623, 
    2648, _, _, 3502, 8232, 3942, 3162, 415, 5960, 8896, 1235, 285, 1730, 
    879, 951, 1436, 601, 648, 2439, 1526, 1013, 287, 366, 1155, 14378, 237, 
    449, 5391, 4125, 689, 1287, 8574, 3211, 58439, 2179, 9821, 6669, 2093, 
    2984, _, 4622, 3541, 7696, 10438, _, 8661, 2776, _, _, _, _, 2706, _, _, 
    2971, _, _, 11804, _, _, 2093, _, 2678, _, _, _, _, _, 1333, 1977, _, 
    877, _, _, _, 316, 453, 489, 5204, 2245, _, 5539, 4526, 7632, 8480, 4439, 
    5062, _, _, 16914, _, _, _, _, 12086, 10476, _, 6169, 5217, _, 3376, 
    2760, _, 27778, 4720, 3102, 660, 783, 21129, 4114, 4390, 3524, 4455, _, 
    _, 4543, 5138, _, _, 6376, 10392, 130287, 112875, 90614, 1991, 1725, 
    3021, 1632, 1327, _, _, _, 2857, 1173, 627, 3423, 1367, 2808, 2398, 1212, 
    2728, 461, 1017, 1029, 258, 2067, 2771, 2755, 1690, 1403, 16664, 2292, 
    2461, 966, 4021, 2976, 3432, _, _, 2798, 2863, _, _, 28948, 8854, 2242, 
    101476, 383, _, 4157, 4735, _, 35231, _, _, _, 681, 742, 1308, 9621, 
    21088, 6649, 254, 593, 4172, 3391, 6303, 8420, 620, 513, 3522, 5883, 
    2830, 5480, 18121, _, 3535, _, 4198, 68538, _, _, _, 6845, _, 980, _, _, 
    788, 1473, 6553, _, 522, _, 860, _, _, _, _, _, _, _, 24873, _, 586, _, 
    1651, 1588, 1229, 1182, 3296, 2294, 4905, 4564, 161957, 522952, 298256, 
    14293, 7466, 8569, 2308, 9165, _, 3619, 5177, 2633, 4058, _, 3742, 54187, 
    _, 1326, 1628, 2055, 31239, _, _, _, _, _, _, _, _, _, _, 318, 1854, 
    1579, 987, 19083, 3836, 432, 452, 373, 417, 453, 256, 589, 649, 1919, 
    926, 1346, 7453, 933, 1322, 1552, 1494, 487, 1874, 4012, _, _, 20344, 
    4280, 1004, _, 11600, 2457, 4943, _, 2746, _, _, _, 3215, 7066, _, _, 
    3617, 46390, _, 1456, 297, _, 1258, 2805, 1593, 553, 801, 37190, 3704, 
    788, 1467, 566, 1289, 2521, 2035, 263, 1066, 4683, 452, 389, _, 640, 
    2871, 355, 1746, 6725, 870, 820, _, 748, 427, 4957, 2006, 1346, 2215, 
    2868, 7797, _, 9621, 10852, 5890, _, _, 2446, _, _, _, _, _, _, _, _, 
    35613, 601, 577, 1146, _, _, 1606, 1100, 1093, 2242, 2788, 2479, 4218, 
    482, 3633, 3295, 3241, _, 1172, 1557, 2706, _, _, 4457, _, _, 5791, 5483, 
    3411, 2363, 1420, 2155, 2291, _, _, _, _, _, _, _, _, 10349, _, _, _, 
    17542, 2693, 2336, 1209, 1503, 7056, 2776, 958, 907, 1433, 725, 1026, 
    4025, 1739, 5884, 1700, 11929, 1292, 405, 1398, _, 4435, 1352, 651, 
    24664, _, 6614, _, 24482, 652, 685, 3392, 12265, 8204, 124541, 3440, 
    3193, _, 1239, _, 1614, 405, 4314, 7113, 4810, 1399, 23749, 808, 8831, 
    9652, 3109, 1822, 4178, 2065, 617, 24399, 24995, 335, 905, 393, 1367, 
    639, 2217, 21280, 10251, 716, 1552, 1626, 3579, _, 1762, 1702, 2080, _, 
    _, _, _, _, _, _, 5284, 5993, 2445, _, 4670, 5204, 17913, 19617, 4747, 
    4473, 4567, 1840, 627, 1934, 4140, 694, 4201, 21729, 8844, 6154, 5714, 
    10538, 4973, 5698, 100647, 5421, 4690, 5506, 94505, 5999, 704, 523, 4114, 
    4428, _, _, 4880, 5420, 80728, 769, 759, 1522, 5717, 300, 315, 1256, 
    1175, 2267, 9452, 1901, 56057, 97484, 2858, 10288, _, 10449, 6415, 469, 
    999, 2235, _, _, _, _, 31760, _, _, _, 1279, 7019, 1382, _, 1890, 811, 
    587, 1420, 1175, 1022, 1477, _, 4034, 20844, 506, _, 685, 5853, 2775, 
    2866, 32778, 7371, 7457, 7527, 473, 8273, 6060, 2630, 1145, 739, 734, _, 
    _, 6432, 1436, 13104, 2992, 2745, _, 26219, 5866, 1784, 9423, 3801, _, _, 
    _, _, _, 4753, _, _, 1128, 406, 759, 1035, 615, _, _, _, 9202, 1925, 
    1359, _, _, 11336, 10083, 6278, 10748, 5926, 3047, 5532, 3985, 8789, 
    1766, 2165, 2092, 2227, 15868, 4939, _, 6393, _, 6447, _, 35327, 3665, 
    2253, 3297, 2050, _, _, 2029, _, _, _, _, _, _, 896, 1163, 1043, 698, 
    937, 892, 1086, 5398, 575, 1281, 465, _, _, 11334, 752, 2891, 2571, 
    10867, 3109, 34280, _, 19627, 11979, 1628, 2915, _, _, _, _, 1623, 4514, 
    _, 57419, 13063, _, 651, _, _, _, _, 16609, 46670, _, _, 29928, _, 
    123353, _, _, 9925, 606, 4778, _, 2612, _, 10516, 2366, _, 3623, 4245, 
    4355, 3443, 3572, 2568, 2671, 4123, 1948, 2162, _, 14252, 10953, 3160, _, 
    736, 650, 321, 1897, 708, 11967, 562, 671, 652, _, 468, 710, 7865, 8652, 
    49999, 8210, _, 12196, 2481, 3700, 22313, 2376, _, _, 11046, _, _, 1983, 
    311, 760, 2804, _, _, _, _, 490, _, _, 3367, 2431, 7758, 6158, 2601, 
    3579, 2798, 1630, _, 8148, 1359, 2118, 1676, 45360, 4203, 11136, _, 
    18936, _, 4069, 2279, 2613, 4262, 8376, _, 7895, 46720, 6870, _, 5631, 
    48146, 15304, 4827, 3753, _, _, 32254, 4414, 5409, 2695, 3195, 1697, 
    2138, 2282, 20459, 1139, 30994, _, 1738, 1757, 2049, 4652, 1955, 7827, 
    1980, 4696, _, 31753, _, _, _, 1351, 385, 321, 1125, 525, 19395, 4735, 
    60830, 6200, 5545, _, 3265, 544, _, 336, _, _, _, 658, _, 1079, _, 1069, 
    2428, 6323, 3691, 2433, _, _, _, _, _, _, _, 13096, 2679, _, _, 7459, 
    6700, 6218, 591, 542, 3222, 4250, 2134, 4789, 7167, 5626, 3794, 24634, 
    4307, 1585, 404, 350, 2325, 2446, 3043, 19275, 972, _, _, _, _, 25367, 
    15069, 37982, 7201, 11496, 17639, _, 2148, _, 141023, 6197, _, 1231, 
    1063, 24938, 11500, 971, _, 2222, _, _, _, _, _, _, _, 3383, _, _, 710, 
    20265, _, 8786, 5079, 1544, 611, 5980, 11530, 4130, 1473, 2413, 527, 974, 
    3804, 31056, 2227, 1774, 1747, _, _, _, _, _, _, 18476, _, 2573, 928, 
    11079, 1800, 364, 2301, _, 414, 2016, 1495, 1961, _, 5672, 19067, 9237, 
    _, 3062, 9754, 2281, 5606, 2457, 2515, 2413, 7956, 341, 1710, 1344, 7913, 
    1910, 10240, 5457, 5538, 6154, 3128, 6744, _, 8316, 625, _, _, _, 11166, 
    _, 16576, 494, 1140, 202, 4556, 9173, 4607, 2057, _, 6242, 2877, 8086, _, 
    2669, _, 45760, _, 1456, _, _, 584, _, 960, _, 1062, 10630, _, 271, 355, 
    1023, 1957, 1924, 1264, 906, 2987, 5122, 1989, 1203, 2994, 4184, 2800, 
    78559, 12292, 5215, 432, 784, 1973, 2133, 4138, 581, 7325, 351, 1509, 
    2460, 532, 2156, 983, 1611, 1759, 2839, 6788, 262, 3962, 1056, 1380, 554, 
    1700, 926, 892, 9751, 22743, 1299, 2737, 5167, 761 ;

 semi_minor_axis = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, 65, 164, 133, 40, 129, 36, 98, 38, 597, _, _, _, _, _, _, _, 1052, _, 
    _, 1001, _, 157, _, _, 41, 89, 192, 21, _, 215, 615, _, 482, _, 507, 61, 
    317, _, _, 873, _, _, 1168, _, _, 1758, _, 1472, 48, 25, 68, 383, 379, 
    25, 235, 222, _, _, _, 431, _, 1507, _, 1158, 500, 399, 646, 46, 456, 99, 
    304, 608, 3439, 146, 1324, 296, 35, 841, 340, 432, 458, 256, 827, 138, 
    53, 533, 588, 209, 619, 724, 159, 181, 187, 26, _, 342, 137, 64, 80, 
    1002, 1064, 211, 170, 3525, 201, _, 182, 55, 79, 163, 600, _, _, _, _, _, 
    _, _, _, _, _, _, 112, 157, 575, 500, _, 922, 150, 187, 27, 4993, 552, _, 
    1553, 1789, 1190, 31, 510, 95, 52, 174, 466, 128, 189, 90, 51, 106, 2890, 
    _, _, _, _, _, _, _, _, _, _, 54, _, _, _, 633, 19, 322, 487, 548, 637, 
    717, 46, 53, 172, 315, 100, 223, 534, 782, 126, 365, _, _, 810, _, _, _, 
    2417, 1914, 331, 627, 192, 1424, 52, 1115, 848, 100, 138, 1223, 125, 64, 
    175, 231, _, 714, 59, 766, 81, 116, 128, 411, 614, _, _, _, _, _, _, _, 
    _, _, _, 4322, 140, 495, _, _, 65, _, 1144, 144, 633, 92, _, 412, 116, _, 
    296, _, 1265, _, 63, 47, 851, 36, 450, 41, 29, 59, 267, 24, 124, _, _, 
    1372, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    4138, _, 244, 2007, 1525, 65, 129, _, 601, 34, 52, 122, 50, 60, 440, 61, 
    192, 553, 1333, 188, 702, _, 139, 166, _, _, _, _, _, _, _, _, _, _, 206, 
    27, 154, 522, 104, 98, 464, 75, 237, 470, 66, 47, 110, 85, 73, 45, 55, 
    49, 628, 33, 39, 329, 60, 193, 176, 160, 43, 120, 598, 595, 507, 161, 
    162, 375, 40, 100, _, 363, _, _, 41, 170, 46, _, 90, _, 49, 200, 324, 
    1006, 40, 211, _, 57, _, 117, _, 76, _, 54, 477, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, 2780, 86, _, _, _, 439, 258, _, _, _, _, 793, _, 
    169, 39, _, 304, 309, _, 244, 34, _, 370, 324, 347, 471, 1419, 662, _, 
    90, 582, 52, _, 807, 913, 2046, _, _, _, _, _, _, _, 1035, _, 145, _, 
    757, 25, 73, 61, 25, 230, 221, 443, 58, 26, _, _, _, _, 553, _, _, 151, 
    _, 928, _, 1990, _, 3647, 381, 163, 1641, 376, 129, _, 173, 182, 217, 86, 
    118, 557, 113, 195, 79, 764, _, _, 1113, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, 68, 987, _, 109, _, 243, _, 71, 
    49, _, 810, 679, 65, 37, 213, 409, 94, _, _, _, 102, 470, _, _, 74, _, 
    90, _, 177, 316, 316, 361, _, _, _, _, _, _, _, _, _, _, _, _, 260, 177, 
    37, 309, _, 386, 24, _, 89, 389, 95, 51, 299, 612, 17, 27, 52, _, _, 638, 
    109, 216, 581, 85, 128, 32, 86, 235, _, 89, 555, 509, 479, 1181, 29, 24, 
    151, 18, 87, 497, 508, 365, 2289, 2334, 1987, 1979, _, _, _, 49, 448, _, 
    109, 618, 790, 85, 527, 223, 437, _, 24, 138, 77, 276, 21, 715, 20, 337, 
    56, 62, 73, _, 540, 798, 464, _, _, _, _, _, _, _, _, 140, _, _, _, _, _, 
    889, _, _, _, 143, _, 351, 316, _, _, _, 585, 29, 116, 88, _, 60, 590, _, 
    628, 418, _, 2755, _, 2380, 158, _, _, _, _, 250, 549, _, 2847, _, 315, 
    _, _, _, _, 167, _, 719, _, _, _, _, 332, 61, 263, 1712, 381, 131, 59, 
    28, 240, 133, 62, 298, 102, 387, 32, 87, 283, 21, 40, 57, 68, 354, 964, 
    117, _, _, _, _, _, _, _, _, _, _, 2356, 276, 60, _, _, 712, _, 780, 174, 
    74, 2135, 142, 67, 56, 105, 57, 61, 657, 43, 807, 66, 50, 98, 526, 448, 
    _, _, _, _, _, _, _, 910, 647, 3157, 46, 442, 438, 207, 369, 136, 51, 30, 
    51, 136, 81, 48, _, 125, 180, _, _, _, _, 134, 242, _, 886, _, 200, 1198, 
    69, 244, 579, 304, 87, 384, 408, 70, 36, 640, 108, 37, 1643, 371, 554, _, 
    _, 230, _, _, 3581, 658, 260, 459, 189, 200, 31, 41, 266, 268, 845, 38, 
    383, 765, 45, 939, 24, 113, _, _, _, _, 388, 3294, 1994, 333, 323, 530, 
    582, _, _, 54, 194, 191, _, 195, _, _, 61, 743, 151, 189, _, 346, 135, _, 
    327, 600, _, 85, 385, 320, 84, 67, 301, 53, 137, _, _, 3269, 60, 356, 
    467, 190, 113, _, 113, 597, 483, 63, 331, 803, 788, 43, 35, 421, 1083, 
    324, 1248, 903, _, _, 916, _, _, _, _, _, _, _, 1326, _, 661, 90, 840, _, 
    88, 189, 1119, 85, 270, 97, 198, _, 220, 193, 72, 109, 28, 112, 93, 326, 
    37, 99, 267, 1435, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 125, 19, 
    218, 130, 986, 384, 38, 190, 18, 136, 98, 75, 127, 196, 18, 42, 77, 92, 
    75, 206, 160, 78, 99, 1264, 1280, 402, 507, _, _, _, _, _, _, _, _, 29, 
    415, _, _, _, _, 28, 71, 245, 248, 32, 224, 18, 19, 17, 338, 480, 98, 
    459, _, 650, _, 870, _, _, 1056, 27, 312, 309, _, 491, _, 166, 138, 162, 
    83, 41, 154, 64, 498, 108, 585, 153, 318, 267, 100, 358, 377, _, 255, 
    368, _, _, 349, 1001, 167, 133, 1072, 772, 308, 95, 208, 165, 271, 203, 
    38, 957, 475, 58, 70, 125, _, 415, _, 106, _, 37, _, 47, _, 273, 690, _, 
    _, _, _, _, 4367, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, 184, _, 1034, _, _, 38, 330, 359, _, _, 193, 184, 
    41, 82, _, 161, 97, _, _, 28, 56, _, _, 197, _, 135, _, 53, 98, _, 160, 
    _, 22, _, 31, _, 37, _, 215, 251, 494, 293, 252, _, _, _, _, _, _, _, 
    2547, 1499, 1487, 51, 379, 208, 705, 57, 275, 181, 184, 65, _, 1002, 144, 
    1741, 47, 91, 69, 330, 166, _, 141, _, 444, 438, 518, 624, 366, _, _, 
    961, _, _, 1134, 1195, 1649, 556, 1837, _, 81, 187, _, 244, 1883, _, 40, 
    _, 60, _, _, _, _, 1131, _, _, _, _, 223, 1086, 157, 186, 4077, 73, 220, 
    45, 464, 59, 65, 114, 1726, 36, 86, _, 443, _, _, 62, _, 1233, _, _, _, 
    _, _, 2755, 43, 305, _, _, _, _, _, _, 145, 996, 150, _, 21, _, 89, _, _, 
    _, 55, 71, 64, 122, 36, 76, 67, 45, 43, 35, _, 111, 24, 478, 60, 90, 173, 
    _, _, 1322, _, _, _, 76, _, _, 30, 75, 115, 271, 274, 83, 18, 241, 823, 
    16, 54, 43, 306, 64, 159, 69, 44, 82, 84, 120, 1661, 404, 348, _, 1732, 
    1160, _, 2125, 262, 40, 22, 485, _, 98, _, _, 370, 529, 623, 840, _, _, 
    _, _, _, 964, 458, _, _, _, _, 286, _, _, 1278, _, _, _, 47, 517, _, 419, 
    _, 732, 50, 108, 83, 31, 33, 47, _, 537, 87, _, _, 132, _, 388, _, 378, 
    _, _, _, _, _, 792, _, 267, _, _, 66, 381, _, _, 206, 168, 100, 99, 70, 
    516, 139, 253, 189, 769, 357, 190, 112, 69, 70, 521, 114, 323, 199, 368, 
    322, _, 19, 71, 133, 32, 30, 44, 26, 14, 62, 188, 617, 808, _, 1151, 92, 
    49, 108, 277, 443, 772, 24, 585, 442, _, 5812, 7242, 5527, _, _, _, 107, 
    433, _, 123, 417, 313, 35, 528, 121, 925, 92, 217, _, _, 221, 296, _, 25, 
    31, 886, _, _, 1131, 1084, 220, _, 4290, 100, 403, _, 1016, _, 684, 843, 
    714, 38, 34, 372, 49, 1919, 227, 102, 449, 937, _, 281, 136, 282, 44, 
    196, 45, 206, 130, 102, 224, 231, 42, 1140, 41, 79, 201, 466, 302, _, _, 
    _, _, _, _, 87, _, _, _, _, 40, 77, 298, 93, 63, 25, 69, _, _, 26, 121, 
    24, 103, 26, 53, 38, 433, 384, 1220, _, _, _, 362, _, _, _, _, _, _, _, 
    _, _, _, _, _, 98, 1045, _, 1961, 24, 278, 127, 528, 1291, 1839, 52, 32, 
    274, 34, 256, 63, 45, 16, 27, 88, 152, _, _, 984, 1220, 848, 842, 9353, 
    348, 905, 1291, 494, 542, 320, 214, 83, 19, 205, 46, 145, 560, _, _, _, 
    _, _, _, 1039, _, 92, 1531, 477, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    1320, 99, 359, 253, _, 60, 62, 800, 1179, 2055, 588, 77, _, 153, 390, _, 
    95, _, 507, 55, _, 113, 273, _, _, 40, 77, _, 98, 195, 627, _, _, _, 976, 
    558, 598, 619, 584, _, 33, 589, _, 409, 442, 520, _, _, _, 113, 211, 553, 
    39, 300, 821, 248, 63, 207, 291, 380, 171, 21, 45, 81, 84, 25, 66, 234, 
    79, 136, 68, 136, _, 6681, _, _, _, _, 92, _, _, 177, _, 35, 188, 292, 
    336, 50, 55, 85, 34, _, 285, 41, 264, 23, 313, 35, _, _, 180, 121, _, 
    314, _, _, 2240, 264, 549, 76, 422, 576, _, _, _, _, _, 2627, 66, 866, 
    635, 64, 213, 149, 264, 65, 29, 110, 948, 602, 29, 27, 34, 243, _, 1952, 
    155, 1095, 3077, 334, 910, 471, _, _, _, _, _, _, _, _, _, _, 698, 995, 
    109, _, 324, _, 114, 438, 349, 1205, 399, 107, 102, _, 462, 240, 1911, 
    561, 880, 66, 125, 53, _, 174, 210, 126, 122, 96, 701, _, _, _, 603, _, 
    802, 3206, 1379, 27, 360, 609, 589, 676, _, 88, _, _, _, _, 1086, 964, 
    739, _, _, _, _, _, 155, 362, _, 1283, _, 95, 35, 282, _, 407, 221, 79, 
    21, 94, 39, 175, 146, _, 465, 148, 135, 55, 319, 1089, 428, 505, _, 126, 
    608, 108, _, 477, 111, 28, 61, 113, 93, 303, 31, 256, 168, 60, 31, 325, 
    761, 1065, 24, 83, 349, 145, _, _, 2985, 80, 90, 72, _, 455, 73, 95, 521, 
    64, 47, 141, 144, 229, 101, 107, 297, 104, 31, 42, 88, 239, 809, 232, _, 
    _, _, 659, _, 2445, 1015, 79, 85, _, 633, 527, 174, 50, _, _, 426, 45, _, 
    846, 59, 869, 135, 204, 105, _, 1123, _, 48, _, 81, _, 21, 83, 169, 351, 
    43, _, _, _, _, _, _, 436, _, 89, _, 211, 216, _, _, 83, _, 45, 152, 176, 
    177, _, 60, 423, 20, 346, 520, 98, _, 310, _, _, 329, 632, 103, 367, 139, 
    81, 1008, 556, 639, 16, 46, 48, 158, _, _, _, _, _, _, _, _, _, _, _, 
    1635, 104, _, 134, 1563, _, 22, 164, 50, _, _, _, _, _, _, _, _, _, _, 
    113, _, _, 549, _, 74, 400, _, 480, _, 499, _, 602, 642, 98, _, 78, _, 
    52, _, 287, _, _, 32, 32, 37, 51, 32, 72, 99, 575, _, 86, _, _, 161, 149, 
    107, 352, 147, _, 225, _, 66, 152, 468, 59, 298, 55, 160, 853, 309, 33, 
    105, 143, 563, 1692, 277, 105, _, _, 1016, 129, 269, 1101, 91, 305, 558, 
    237, _, 626, 459, _, 70, 63, 291, 106, 474, 589, 194, 78, 51, _, 49, 37, 
    _, 461, 590, 696, _, 1147, 207, _, _, _, _, 907, _, 52, _, 523, _, 1743, 
    3089, 37, 196, 550, _, 592, 102, 73, 178, 309, 50, 124, 87, 57, 114, 104, 
    1119, 48, 462, 1077, _, _, _, _, _, 129, _, 521, 78, 678, 184, _, _, _, 
    _, _, _, _, 1573, 1846, 1759, 246, 444, 100, 1982, 169, _, 1201, 47, 22, 
    131, 42, 800, 62, 53, 1019, 27, _, _, 463, 288, 746, _, _, _, _, _, 77, 
    718, 65, 29, _, 297, 355, 70, 119, 221, 306, 990, 233, 173, 95, 158, 319, 
    _, _, 204, 46, 41, 200, 1401, 604, 106, 108, 96, _, _, _, _, _, _, 47, 
    934, 75, 65, 394, 143, 333, 112, 688, 62, 692, 46, 102, 164, _, 538, _, 
    585, _, 84, _, _, _, _, _, _, _, _, 1005, 887, 2409, 1097, _, _, _, 3564, 
    2188, 122, 1900, 3177, 2817, _, _, _, _, 27, 21, 64, _, 28, 92, 48, _, _, 
    86, 1113, 4147, 3780, _, 48, 83, 114, _, 15, 1034, _, _, 2289, 46, 1261, 
    984, 25, _, _, _, _, 58, 764, _, 23, 283, 307, 382, 424, _, 659, 472, 
    475, 116, 597, 852, 66, 86, 33, 262, 60, 50, 56, 33, _, 83, 98, _, _, _, 
    982, _, _, _, 1161, _, 918, _, 178, _, _, _, _, 111, 225, _, 195, _, 
    1621, _, _, 367, _, 78, 244, _, 143, 594, _, 650, 671, 645, 227, _, _, 
    60, _, 335, 1163, 1634, 1091, 228, 406, 431, 58, 514, 980, 1669, 67, _, 
    65, _, 224, 248, 83, _, _, 1491, 918, _, 591, 625, _, _, _, 845, 893, 
    928, 47, 35, _, _, _, _, _, _, 1918, 1591, 126, 72, 464, 650, 375, 172, 
    109, 178, 117, 91, 145, 722, 115, 461, 378, _, 85, 103, 74, 107, 43, 59, 
    852, 131, _, _, _, 1470, 65, 798, 65, 69, 381, 637, _, _, 132, 39, 98, 
    227, 71, 55, 41, 66, 47, 34, 30, 272, 85, _, _, 19, 204, _, 1077, 22, _, 
    20, 139, _, 127, 72, 431, 25, 30, 221, 771, 767, _, 1213, _, _, _, 979, 
    1053, 278, 2265, 3036, 311, _, 489, 929, 614, 622, 29, 490, 95, _, 63, 
    265, 228, _, 994, 114, 219, 69, _, 122, 69, 62, _, 83, 285, 1863, 1185, 
    _, _, _, _, 917, 1576, _, _, _, 1048, _, _, 583, 1170, 65, 36, _, _, _, 
    83, _, _, 557, _, 707, 801, _, 827, _, _, 54, _, _, 218, 120, _, 154, 
    453, _, 1528, 838, _, 853, 147, 250, 419, 218, _, 6137, _, 56, 402, _, 
    131, 360, 736, 22, 111, 151, 220, 49, 87, 117, 148, _, 201, 108, _, 86, 
    90, 426, _, 506, _, 421, _, _, _, _, _, _, _, 2063, 181, 53, _, _, _, _, 
    118, 494, 916, 1676, 604, _, 331, _, 203, 225, 112, 267, 89, 262, 63, 
    345, 40, 88, 311, 28, 79, 42, 229, 223, 960, _, _, _, _, _, _, _, 56, 
    134, 78, 85, 418, 39, 85, _, 44, 61, _, _, 106, 174, 21, _, 93, 159, 
    2375, 131, 771, _, _, _, _, _, _, _, _, _, _, _, _, 3062, _, _, 97, 772, 
    1234, 1633, 427, 396, 448, 487, 426, 160, 531, 142, 31, 37, 32, 360, 23, 
    166, 137, 138, 594, 829, 162, 116, 166, 1985, 156, 398, 91, 98, 79, 69, 
    191, 190, 812, 107, 504, 298, 87, 102, 60, 68, 30, 686, 107, 133, 118, 
    115, _, _, _, _, _, _, _, _, _, _, 693, 93, 406, 68, 108, 882, 953, _, 
    1376, 21, 229, 934, 70, 128, 56, 487, 229, 51, 65, 32, _, 55, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, 2616, 2892, _, _, 1958, _, _, 1614, 128, 247, 
    238, 969, 579, 58, 295, 55, 67, 447, 100, 97, 125, 270, 190, 396, 163, 
    55, 64, 165, 153, _, 215, 1204, _, _, _, _, _, _, 1832, _, 321, _, 126, 
    65, 18, 106, _, 198, 626, _, 385, 490, _, 74, _, 40, _, 243, _, 392, 306, 
    289, _, 4397, 3346, 3698, 4159, 560, 556, _, _, _, _, _, 105, _, _, 591, 
    157, _, _, 508, 55, 157, 76, 47, 266, 42, 45, 245, 676, 599, 658, 47, _, 
    _, _, _, _, _, _, 201, 730, _, _, 45, 105, 25, 176, 69, 248, _, 239, 
    1418, 517, 80, 21, _, 286, _, 373, _, _, 208, 543, _, 1363, 121, _, _, _, 
    _, 2504, 184, 304, 43, 450, 368, 65, 164, 96, 45, 79, 29, 40, 75, 90, 19, 
    278, 25, 41, 36, 45, 439, 225, 202, 654, _, _, _, 17, _, 186, _, 525, 
    652, 1472, 223, 170, 45, 265, _, 1041, 47, 76, 55, 302, 59, _, 81, 89, 
    103, 171, 343, 449, 563, 680, _, _, _, _, _, _, _, _, _, _, 510, 108, _, 
    112, 116, 804, 366, _, 89, 340, _, 1554, 794, 16, 99, 129, 41, 28, 144, 
    _, 766, 107, _, 224, 234, _, _, _, _, _, _, _, _, _, 1548, 266, 1958, 
    108, _, 32, _, 237, _, 126, 152, 452, _, 30, 274, 351, _, 141, 22, 288, 
    38, 105, 22, 50, 75, _, 56, _, 79, 98, 384, 318, 2232, _, 2339, _, _, _, 
    _, _, 781, _, 238, _, _, _, _, _, _, _, _, _, 219, 214, 48, 506, 638, 76, 
    _, 62, _, _, 77, 441, 200, 27, _, _, 79, 99, _, 120, 205, _, _, 348, _, 
    642, 609, 68, 438, 153, 427, 631, _, _, 251, 1451, 575, 2153, 1467, 275, 
    559, 62, 459, _, 929, _, _, 1122, 261, 57, 74, 53, 152, 35, 75, 321, 83, 
    47, 1063, 131, 257, 1207, _, 2405, _, 492, 335, _, _, _, 614, 812, 800, 
    100, 474, 161, 80, 444, 806, 75, 615, 828, 715, 658, 77, 188, 291, 47, 
    147, _, 627, 642, 79, 480, 817, _, _, _, _, _, _, _, _, 229, 299, _, 705, 
    _, _, _, 96, 511, 265, 284, _, 424, 511, 96, 102, 151, 335, 83, 237, 40, 
    269, 22, 365, 367, _, _, 491, 85, 1189, 100, _, 1239, 1060, _, _, 984, 
    28, 190, 1167, 439, 705, 741, 186, 1400, 101, _, 32, 369, 111, 588, 103, 
    56, 192, 22, 30, 31, 214, 42, 1032, 810, 104, 176, 114, _, _, _, _, _, _, 
    944, 67, 171, _, _, 143, 118, _, _, 78, 114, 179, 69, _, 57, _, _, 167, 
    _, 277, 154, _, 219, 73, _, 377, _, 89, 588, _, _, _, _, _, _, _, _, _, 
    286, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 1777, 83, _, _, 62, _, 
    1429, _, 23, 88, 466, 977, 881, 530, 544, 314, 59, 57, 83, 783, 620, _, 
    1480, 162, 25, 349, 108, _, 132, _, _, 56, _, 76, 853, 95, 302, 248, 157, 
    98, 198, 106, 30, _, 51, 21, 93, 114, _, _, 231, 834, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, 97, _, _, 364, 882, 36, 228, 416, 533, 537, 
    464, 461, 572, 41, 45, 368, 155, 209, 644, 29, 195, _, 195, _, _, _, _, 
    165, 1292, 114, 171, 32, 139, 83, 815, _, 393, 251, 61, 112, _, _, 54, 
    136, 73, _, 89, _, _, 468, 48, 235, 398, 91, 58, 92, _, 292, _, _, 109, 
    231, _, _, 274, _, 3118, 201, 311, 191, 35, 52, 60, 131, 199, 211, 62, 
    39, 28, 108, 793, 54, _, 284, 982, 1905, _, 2386, 2210, 189, 105, 90, 65, 
    897, 742, 622, 25, _, _, 370, _, 433, 491, _, 529, 84, 91, _, 448, _, 
    565, 586, 646, 135, 382, 361, 539, 387, 44, 51, 82, 63, 268, 460, 1176, 
    84, 16, 189, 294, 103, 101, 71, 63, 36, 532, 160, 632, _, _, 86, 22, 414, 
    172, 71, 403, _, _, _, 802, 32, 42, 134, 105, 585, 1990, 1900, 6602, 
    4288, 3834, 30, 42, 76, 115, 484, 26, _, 123, 27, 48, 206, 100, 130, 293, 
    42, 706, 506, 529, _, 59, _, _, _, 3504, 120, 324, 947, _, 40, _, 42, _, 
    79, 105, 69, _, 173, 178, 1898, 488, 142, 485, 120, 93, 81, _, _, _, 
    1177, _, _, 38, _, _, _, _, 558, 18, 159, 43, _, 49, 482, 74, 39, 130, _, 
    _, 702, 69, 92, 84, 1849, 147, 452, 2058, _, 5375, 468, 67, 76, 82, 210, 
    2430, 2557, 20, 67, 264, 481, 457, 610, 514, 334, 43, 600, 579, 537, _, 
    _, _, _, 154, 121, 507, 76, 52, 69, _, _, _, _, 1645, 314, 334, 506, 140, 
    344, 1398, 111, 83, 103, 160, _, 73, 238, 28, 130, 143, 61, 71, 53, 38, 
    _, 227, 64, 352, _, 164, _, 175, 258, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, 1353, _, _, _, 28, _, 336, _, 280, 226, _, 235, 132, 1387, 43, 564, 
    79, 20, 107, 510, 100, 357, 47, 46, 149, 88, 37, 403, 138, 230, 416, _, 
    _, _, _, 8547, _, 219, _, 990, 549, 90, 240, 124, 70, 76, 264, 896, 50, 
    35, 33, 133, 116, 201, 27, 70, 376, 236, 98, 200, _, _, _, _, _, _, _, _, 
    51, _, 21, _, 147, 353, _, _, 341, 333, 212, _, _, 36, 112, _, 27, _, 
    353, 61, 53, _, 379, _, 39, 70, 205, 696, 907, _, 312, _, 2226, _, _, 
    398, 512, 523, _, _, 24, _, _, 340, 829, _, 35, _, _, 72, 69, _, _, 164, 
    40, 59, _, 255, _, _, 108, 2929, 2475, 131, 373, _, _, _, 705, 1057, _, 
    84, 1249, _, 86, 80, 137, 55, _, 33, _, _, _, 76, 38, _, 262, 76, 141, 
    3470, _, 425, 409, _, _, _, 1085, 547, _, _, 811, _, _, 27, _, 239, _, 
    111, _, 114, 56, 139, 505, 24, 102, 351, 835, 1475, 1123, 160, 449, _, _, 
    _, _, 2921, 2533, _, 811, 1057, 184, _, 969, _, 21, _, 50, 118, 2217, 
    192, 752, 582, 97, 34, 369, 64, _, 383, 605, _, _, _, 148, _, _, 986, 
    103, 107, 214, 185, _, _, _, _, _, _, 134, _, 194, 429, 814, _, _, 30, 
    134, 133, 66, 420, 504, 451, 60, 51, _, 28, _, 246, _, _, 624, _, _, 81, 
    174, 627, 62, _, 573, 455, 46, 175, 68, 296, _, 200, 34, _, _, _, _, _, 
    946, _, 138, _, 86, 37, 58, 632, 1280, 41, 43, 59, 347, 24, _, 1281, 910, 
    _, 269, 1931, 1559, 2562, 1953, 26, 2838, 259, 75, 179, 109, 234, 172, 
    415, 1106, 181, 421, 36, 49, 70, 41, 216, 40, _, 437, 378, 47, 60, 467, 
    800, 225, _, _, _, _, 926, _, _, 683, 443, 882, 139, 156, 228, 100, 128, 
    _, _, _, _, 125, 1112, _, 76, 96, 220, 77, 149, 434, 323, 27, 230, 426, 
    241, 30, 30, 36, 83, 153, 91, 343, 67, 147, 206, 47, 101, 25, 91, 238, 
    173, 1915, 1667, _, 63, 259, 311, 40, 121, _, 171, 47, 302, 64, 236, 506, 
    71, 85, 476, 168, 915, 44, 346, 599, 72, _, 587, 117, _, 245, 147, _, _, 
    1029, 43, 747, 115, 385, 225, 244, 144, _, 100, 62, 34, 28, 615, 54, 64, 
    95, 164, _, 1116, _, _, _, 4503, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, 8075, 7131, _, 68, 623, 618, 120, 304, 375, 128, 628, 23, 74, _, 49, 
    87, _, _, 79, _, 34, _, 151, 755, _, 1454, 98, 337, 42, _, _, 117, _, 
    147, _, _, _, _, 2982, 447, 444, 619, 1133, 1308, 1177, _, 879, _, 30, _, 
    212, 128, 60, 51, 94, _, 176, 92, 101, 2527, 448, 165, _, _, 1327, 59, 
    826, 17, 54, 1556, 1519, 211, 246, 400, 290, 588, 402, 33, 248, 58, 281, 
    574, 79, 42, 129, 16, 145, 91, 46, 277, 45, 34, 30, 704, 1296, 55, 180, 
    1689, 161, 197, _, 43, 90, 1874, 323, _, 89, 192, _, _, _, _, 499, _, _, 
    666, _, _, 165, _, _, 1042, _, 24, _, _, _, _, _, 144, 777, _, 140, _, _, 
    _, 66, 42, 189, 2482, 561, _, 459, 33, 89, 99, 256, 134, _, _, 612, _, _, 
    _, _, 1188, 1033, _, 804, 851, _, 61, 90, _, 47, 251, 252, 114, 291, 23, 
    278, 314, 442, 317, _, _, 518, 873, _, _, 1103, 678, 675, 614, 530, 45, 
    315, 90, 127, 645, _, _, _, 397, 79, 108, 1265, 114, 236, 259, 418, 320, 
    68, 264, 263, 93, 503, 74, 1211, 97, 292, 36, 243, 408, 515, 121, 171, 
    86, _, _, 644, 602, _, _, 72, 112, 532, 34, 68, _, 835, 573, _, 24, _, _, 
    _, 72, 97, 349, 384, 227, 49, 228, 236, 128, 515, 61, 71, 273, 145, 41, 
    1080, 555, 16, 18, _, 551, _, 1104, 54, _, _, _, 412, _, 358, _, _, 161, 
    362, 22, _, 412, _, 183, _, _, _, _, _, _, _, 104, _, 120, _, 206, 216, 
    59, 233, 187, 108, 1177, 956, 63909, 51021, 93980, 94, 126, 28, 292, 58, 
    _, 325, 333, 1201, 1824, _, 1639, 65, _, 230, 718, 696, 75, _, _, _, _, 
    _, _, _, _, _, _, 204, 180, 406, 581, 45, 318, 332, 103, 53, 136, 49, 
    183, 159, 43, 517, 26, 21, 21, 62, 51, 36, 117, 73, 354, 184, _, _, 18, 
    28, 128, _, 24, 256, 99, _, 481, _, _, _, 1024, 551, _, _, 1215, 23, _, 
    32, 64, _, 303, 360, 1022, 74, 190, 74, 232, 59, 369, 47, 78, 113, 348, 
    96, 284, 95, 162, 135, _, 64, 93, 123, 362, 43, 41, 180, _, 65, 207, 154, 
    362, 125, 110, 83, 1736, _, 2346, 2758, 167, _, _, 1214, _, _, _, _, _, 
    _, _, _, 123, 190, 262, 362, _, _, 252, 313, 199, 604, 257, 27, 37, 62, 
    51, 804, 194, _, 829, 386, 90, _, _, 28, _, _, 68, 27, 101, 603, 130, 
    292, 449, _, _, _, _, _, _, _, _, 1560, _, _, _, 53, 929, 271, 390, 259, 
    187, 26, 58, 53, 29, 82, 244, 40, 83, 20, 37, 63, 207, 79, 326, _, 93, 
    59, 115, 89, _, 522, _, 86, 38, 69, 851, 214, 518, 85, 368, 477, _, 24, 
    _, 412, 198, 1118, 294, 64, 224, 1647, 152, 2153, 1988, 123, 243, 1073, 
    261, 372, 52, 234, 193, 191, 37, 87, 54, 542, 35, 35, 39, 390, 373, 219, 
    _, 857, 482, 107, _, _, _, _, _, _, _, 2301, 2028, 175, _, 1147, 1350, 
    840, 88, 990, 1072, 1060, 528, 168, 380, 69, 36, 420, 5712, 16, 180, 65, 
    61, 193, 1047, 42, 188, 539, 802, 105, 1358, 39, 70, 1456, 1861, _, _, 
    1531, 1129, 40, 84, 160, 402, 158, 227, 256, 61, 69, 57, 57, 472, 1616, 
    83, 1121, 1924, _, 2063, 132, 199, 72, 355, _, _, _, _, 4280, _, _, _, 
    834, 61, 228, _, 171, 70, 79, 102, 203, 72, 188, _, 1121, 224, 166, _, 
    129, 56, 466, 806, 354, 3200, 1221, 2558, 96, 343, 48, 47, 149, 62, 62, 
    _, _, 49, 45, 30, 215, 246, _, 29, 144, 25, 69, 456, _, _, _, _, _, 1116, 
    _, _, 43, 217, 173, 96, 147, _, _, _, 423, 138, 295, _, _, 122, 868, 
    1639, 2768, 1370, 251, 770, 1925, 44, 385, 594, 708, 755, 139, 220, _, 
    79, _, 1549, _, 146, 91, 471, 222, 331, _, _, 96, _, _, _, _, _, _, 197, 
    357, 169, 54, 259, 147, 178, 322, 71, 80, 168, _, _, 77, 47, 738, 661, 
    62, 333, 594, _, 1465, 432, 750, 650, _, _, _, _, 367, 1440, _, 147, 100, 
    _, 394, _, _, _, _, 4393, 2484, _, _, 2030, _, 37, _, _, 507, 164, 41, _, 
    89, _, 53, 48, _, 310, 266, 299, 493, 573, 463, 173, 19, 321, 437, _, 50, 
    40, 343, _, 193, 38, 46, 387, 46, 315, 40, 97, 162, _, 86, 51, 36, 33, 
    31, 600, _, 31, 382, 299, 974, 1688, _, _, 3614, _, _, 413, 68, 356, 211, 
    _, _, _, _, 143, _, _, 912, 940, 98, 144, 134, 106, 491, 67, _, 18, 112, 
    103, 114, 68, 39, 2850, _, 3128, _, 33, 458, 572, 460, 1030, _, 1012, 
    302, 60, _, 1002, 29, 85, 390, 406, _, _, 112, 330, 70, 242, 693, 137, 
    656, 779, 85, 442, 121, _, 303, 349, 334, 16, 446, 97, 69, 1261, _, 149, 
    _, _, _, 46, 90, 73, 26, 64, 172, 2393, 107, 360, 96, _, 1379, 78, _, 
    135, _, _, _, 66, _, 139, _, 74, 609, 1405, 295, 776, _, _, _, _, _, _, 
    _, 3831, 174, _, _, 1400, 1104, 67, 39, 68, 258, 129, 223, 459, 1809, 
    1348, 286, 82, 181, 97, 114, 85, 657, 648, 836, 195, 61, _, _, _, _, 290, 
    305, 43, 445, 69, 28, _, 463, _, 21, 1596, _, 433, 690, 37, 64, 62, _, 
    609, _, _, _, _, _, _, _, 576, _, _, 137, 69, _, 626, 66, 36, 156, 1553, 
    49, 139, 205, 41, 122, 69, 955, 64, 90, 419, 434, _, _, _, _, _, _, 75, 
    _, 42, 245, 317, 428, 149, 57, _, 50, 260, 510, 125, _, 1354, 170, 433, 
    _, 1239, 312, 1018, 22, 240, 40, 65, 357, 113, 77, 104, 21, 246, 88, 
    1210, 1211, 1386, 80, 239, _, 67, 187, _, _, _, 205, _, 113, 132, 39, 
    158, 805, 36, 389, 40, _, 31, 468, 102, _, 959, _, 65, _, 101, _, _, 71, 
    _, 241, _, 134, 1144, _, 249, 187, 675, 834, 827, 152, 103, 173, 195, 49, 
    43, 814, 1124, 743, 52, 1045, 260, 112, 68, 480, 606, 1000, 122, 38, 115, 
    847, 781, 97, 648, 30, 411, 413, 389, 191, 136, 72, 22, 326, 64, 125, 
    290, 64, 445, 134, 308, 140, 54, 228 ;

 time = 943887902, 943890596, 943895188, 943916305, 943919046, 943921935, 
    944017178, 944018179, 944053798, 944058772, 944061977, 944062868, 
    944064655, 944075880, 944076834, 944081456, 944082456, 944083536, 
    944100789, 944101675, 944109368, 944111559, 944141661, 944167557, 
    944186635, 944189797, 944191817, 944193898, 944194839, 944195867, 
    944197862, 944206869, 944207758, 944226670, 944305130, 944307911, 
    944309980, 944315969, 944319798, 944320841, 944323703, 944326388, 
    944328175, 944329075, 944359032, 944360185, 944362551, 944365099, 
    944366054, 944366600, 944367283, 944368329, 944391822, 944392048, 
    944392918, 944393937, 944394926, 944395935, 944396819, 944397768, 
    944397769, 944398937, 944401248, 944402906, 944403175, 944403612, 
    944404112, 944405014, 944415439, 944415538, 944415981, 944416096, 
    944416655, 944416893, 944421002, 944421596, 944422300, 944422680, 
    944423367, 944425656, 944429246, 944432877, 944433906, 944435147, 
    944438058, 944440101, 944440106, 944442136, 944444029, 944446050, 
    944455926, 944458085, 944458491, 944458935, 944461109, 944463351, 
    944463351, 944463677, 944464820, 944464820, 944471773, 944480592, 
    944481478, 944482266, 944482376, 944488342, 944493358, 944494241, 
    944494822, 944494822, 944500809, 944500919, 944502437, 944507906, 
    944508703, 944510631, 944512670, 944512747, 944513773, 944514327, 
    944516672, 944518629, 944518853, 944519894, 944520213, 944524478, 
    944525797, 944530379, 944530383, 944531254, 944531720, 944532004, 
    944534541, 944537003, 944537585, 944537585, 944537609, 944542236, 
    944543443, 944544162, 944545997, 944549360, 944551955, 944554179, 
    944555667, 944572551, 944578554, 944579629, 944580560, 944582546, 
    944584678, 944585896, 944586682, 944587481, 944587541, 944588818, 
    944594222, 944595170, 944596984, 944602501, 944606099, 944607900, 
    944612409, 944613307, 944614198, 944615108, 944615311, 944616188, 
    944617139, 944617382, 944617799, 944619413, 944620978, 944621757, 
    944622085, 944623110, 944623374, 944624097, 944625162, 944627437, 
    944627437, 944627906, 944628575, 944628739, 944629124, 944631209, 
    944633142, 944633264, 944634083, 944634773, 944635144, 944637022, 
    944639296, 944642201, 944643171, 944646057, 944647025, 944649258, 
    944652066, 944663418, 944669039, 944669955, 944700613, 944701724, 
    944702456, 944704337, 944705325, 944706291, 944707826, 944712081, 
    944714125, 944715184, 944716657, 944717868, 944718710, 944718710, 
    944719889, 944721053, 944722160, 944724250, 944724550, 944726128, 
    944728659, 944730106, 944730372, 944732165, 944736174, 944736660, 
    944738465, 944739357, 944783995, 944785183, 944787397, 944787483, 
    944790826, 944793250, 944793499, 944794585, 944795556, 944796768, 
    944797095, 944797853, 944799107, 944799606, 944800556, 944801400, 
    944802180, 944802985, 944803306, 944803816, 944805152, 944806724, 
    944807270, 944811141, 944812789, 944845373, 944857730, 944860738, 
    944861637, 944862557, 944863452, 944867277, 944868259, 944869269, 
    944870165, 944872670, 944873344, 944875020, 944878209, 944879112, 
    944879119, 944880006, 944880461, 944880938, 944881502, 944881622, 
    944883699, 944884220, 944885234, 944885515, 944886057, 944886415, 
    944886655, 944887315, 944887476, 944887840, 944889023, 944890251, 
    944891571, 944892026, 944892526, 944893641, 944893846, 944894892, 
    944896341, 944896859, 944898741, 944899563, 944904606, 944921975, 
    944923066, 944924049, 944925289, 944926199, 944927299, 944931991, 
    944932876, 944935555, 944936628, 944937657, 944938590, 944941332, 
    944950074, 944950983, 944951975, 944952838, 944953821, 944954801, 
    944955856, 944959293, 944964583, 944964765, 944966057, 944966057, 
    944966881, 944971027, 944971240, 944972006, 944972729, 944975691, 
    944978015, 944978041, 944978158, 944978910, 944980096, 944981492, 
    944984191, 944984191, 944984242, 944987455, 944989193, 944989853, 
    944989946, 944991121, 944992025, 944994948, 945024499, 945025457, 
    945030394, 945031338, 945032300, 945036159, 945042595, 945044651, 
    945050657, 945051430, 945054661, 945056663, 945056663, 945057118, 
    945057664, 945057846, 945059211, 945060530, 945062669, 945062851, 
    945062851, 945063306, 945063748, 945065308, 945066559, 945068629, 
    945068811, 945069676, 945071223, 945072497, 945075181, 945106756, 
    945106756, 945107199, 945107527, 945112607, 945112607, 945113215, 
    945130413, 945130413, 945130673, 945136437, 945136504, 945138756, 
    945140066, 945140597, 945141524, 945142240, 945142552, 945143434, 
    945143455, 945145640, 945145640, 945147262, 945148121, 945148774, 
    945149949, 945151812, 945153158, 945153480, 945153936, 945154375, 
    945155380, 945156177, 945156356, 945157092, 945157821, 945160343, 
    945165271, 945187564, 945190637, 945192701, 945193627, 945194669, 
    945201629, 945202510, 945204330, 945205316, 945208257, 945211216, 
    945213269, 945214319, 945215338, 945216242, 945216495, 945217326, 
    945218367, 945219333, 945221243, 945221536, 945221995, 945222270, 
    945223140, 945224071, 945225195, 945225809, 945226105, 945227368, 
    945227368, 945227970, 945228169, 945229115, 945229995, 945230846, 
    945231722, 945233040, 945233406, 945233406, 945234261, 945235032, 
    945236875, 945237478, 945238318, 945239018, 945239327, 945241074, 
    945241474, 945241884, 945242990, 945245182, 945254379, 945255299, 
    945257095, 945258017, 945258904, 945259812, 945260702, 945260733, 
    945262516, 945266915, 945270056, 945270695, 945272303, 945272837, 
    945276646, 945277959, 945278855, 945278855, 945280896, 945282739, 
    945282739, 945302941, 945303890, 945304823, 945308461, 945309209, 
    945310256, 945311180, 945312045, 945312061, 945313769, 945314886, 
    945315050, 945315777, 945316572, 945318417, 945318452, 945320056, 
    945320838, 945320861, 945321544, 945322023, 945322173, 945324324, 
    945324393, 945326597, 945326751, 945328041, 945328201, 945330288, 
    945332563, 945332817, 945333714, 945334280, 945334616, 945335516, 
    945338224, 945342714, 945345443, 945350825, 945355340, 945358135, 
    945359035, 945359945, 945361746, 945363536, 945366281, 945367287, 
    945369276, 945371658, 945372712, 945373644, 945374530, 945376377, 
    945377275, 945389820, 945390783, 945393608, 945393608, 945397169, 
    945399536, 945399894, 945400498, 945400974, 945401450, 945401537, 
    945402820, 945403324, 945405670, 945405670, 945406627, 945406769, 
    945407408, 945408940, 945409481, 945409617, 945410597, 945411685, 
    945411818, 945412494, 945412630, 945413536, 945413643, 945414566, 
    945415350, 945415435, 945418460, 945418597, 945419325, 945421645, 
    945446114, 945447902, 945449828, 945450811, 945451675, 945453608, 
    945464243, 945467204, 945468120, 945469071, 945470077, 945475247, 
    945481901, 945485218, 945485341, 945486168, 945486451, 945486729, 
    945487851, 945488335, 945489037, 945491165, 945492287, 945492287, 
    945494570, 945496984, 945498015, 945498362, 945500578, 945501175, 
    945502089, 945502951, 945506985, 945520544, 945523365, 945526277, 
    945529098, 945532556, 945621370, 945622271, 945625053, 945626914, 
    945627237, 945628427, 945629609, 945633097, 945633241, 945633963, 
    945634351, 945635372, 945639166, 945640149, 945640244, 945641445, 
    945645228, 945645978, 945646230, 945647366, 945647574, 945648497, 
    945649514, 945650891, 945653413, 945654436, 945656431, 945657026, 
    945657638, 945660166, 945662600, 945662662, 945663422, 945663714, 
    945663983, 945664911, 945666413, 945667550, 945668688, 945668961, 
    945669552, 945669871, 945671509, 945672146, 945673059, 945674277, 
    945674714, 945675887, 945677042, 945686481, 945687357, 945689162, 
    945690188, 945691075, 945691976, 945693111, 945694955, 945695455, 
    945696900, 945698729, 945699611, 945700505, 945701628, 945701629, 
    945702719, 945703764, 945706228, 945706429, 945707380, 945707380, 
    945707380, 945708536, 945710565, 945711475, 945712589, 945713477, 
    945713734, 945714772, 945716508, 945718505, 945718645, 945719674, 
    945719947, 945720476, 945724112, 945724371, 945725131, 945725942, 
    945726535, 945727441, 945728551, 945729417, 945730337, 945730443, 
    945730547, 945731235, 945731526, 945732114, 945732518, 945733077, 
    945734072, 945734934, 945735834, 945736257, 945736754, 945736904, 
    945738545, 945740337, 945741241, 945742139, 945742189, 945742337, 
    945742550, 945744595, 945745004, 945747839, 945748319, 945748774, 
    945749092, 945750093, 945751003, 945752186, 945753733, 945754416, 
    945755053, 945756024, 945756964, 945758147, 945759853, 945761150, 
    945761969, 945762515, 945764335, 945780169, 945785386, 945786360, 
    945798494, 945799503, 945806045, 945807171, 945808148, 945810011, 
    945810936, 945815110, 945823676, 945827631, 945827965, 945828453, 
    945829331, 945829628, 945832116, 945833113, 945833451, 945833972, 
    945834921, 945835376, 945838971, 945839335, 945840882, 945841200, 
    945841382, 945843839, 945845022, 945845659, 945847069, 945847206, 
    945847297, 945851210, 945853439, 945893858, 945894938, 945895856, 
    945896993, 945900851, 945901768, 945902786, 945912561, 945912585, 
    945914062, 945918298, 945919742, 945920110, 945920580, 945920715, 
    945924198, 945924689, 945925840, 945926615, 945926783, 945930167, 
    945931725, 945932088, 945932548, 945932870, 945934988, 945935969, 
    945936840, 945937788, 945938670, 945938893, 945943446, 945943447, 
    945945503, 945957592, 945960896, 945963646, 945966966, 945967864, 
    945967864, 945969896, 945970213, 945970578, 945973761, 945973785, 
    945976151, 945976251, 945976481, 945979897, 945993681, 945997495, 
    945997997, 945998909, 945999450, 946000691, 946002661, 946003478, 
    946004575, 946005342, 946005933, 946006350, 946009310, 946009384, 
    946010527, 946011527, 946011527, 946013755, 946015328, 946015454, 
    946018265, 946021404, 946039725, 946045382, 946049344, 946053898, 
    946056596, 946057496, 946074019, 946085220, 946086404, 946088144, 
    946088894, 946088894, 946091109, 946092200, 946092722, 946093908, 
    946094311, 946094876, 946094876, 946096991, 946097947, 946098894, 
    946100032, 946100349, 946100349, 946101139, 946103008, 946103386, 
    946104216, 946104975, 946105761, 946106696, 946110438, 946113927, 
    946124111, 946130193, 946135025, 946136236, 946141107, 946141819, 
    946143910, 946144112, 946155511, 946156494, 946168103, 946170905, 
    946173052, 946173495, 946174036, 946176150, 946176609, 946176819, 
    946177859, 946179410, 946179962, 946183198, 946184448, 946185018, 
    946185552, 946185647, 946187808, 946189965, 946191809, 946194143, 
    946195817, 946196282, 946197296, 946197949, 946208099, 946209000, 
    946209995, 946210873, 946214947, 946215866, 946220595, 946220688, 
    946226342, 946226810, 946226974, 946227658, 946228172, 946228686, 
    946256571, 946258102, 946262443, 946263467, 946263969, 946264054, 
    946264325, 946265142, 946267343, 946268554, 946269408, 946269934, 
    946270068, 946270795, 946272887, 946275376, 946275425, 946275889, 
    946275889, 946292865, 946309688, 946315083, 946315981, 946316885, 
    946317803, 946318678, 946321399, 946322301, 946325950, 946332959, 
    946333859, 946334764, 946336555, 946342244, 946348068, 946348568, 
    946348705, 946354392, 946354529, 946354574, 946354938, 946355120, 
    946355939, 946358032, 946360535, 946360671, 946360944, 946361172, 
    946362036, 946363947, 946445117, 946445636, 946445636, 946446646, 
    946447147, 946449623, 946450886, 946451668, 946452893, 946453290, 
    946453663, 946455649, 946456748, 946461059, 946463056, 946464969, 
    946466095, 946472522, 946480226, 946484128, 946484818, 946485900, 
    946486797, 946487839, 946489356, 946489919, 946490574, 946490574, 
    946495238, 946495962, 946497029, 946497150, 946499115, 946501149, 
    946503237, 946504764, 946507118, 946507452, 946508885, 946513460, 
    946513953, 946514408, 946517275, 946518870, 946519634, 946520791, 
    946520791, 946522333, 946522653, 946525467, 946526483, 946526541, 
    946528712, 946529783, 946530557, 946530728, 946532181, 946532486, 
    946534419, 946535756, 946537004, 946538353, 946538780, 946540331, 
    946541438, 946547223, 946550641, 946553117, 946558679, 946577995, 
    946589278, 946599293, 946599995, 946603835, 946605397, 946605824, 
    946607900, 946608005, 946609846, 946611397, 946611697, 946612294, 
    946613504, 946614108, 946615320, 946616351, 946617341, 946618210, 
    946619488, 946620021, 946620072, 946620907, 946621738, 946621799, 
    946623522, 946623598, 946624215, 946624510, 946625788, 946626108, 
    946637913, 946638775, 946639776, 946641930, 946642837, 946643585, 
    946646045, 946647061, 946648038, 946649017, 946650021, 946653719, 
    946654633, 946655581, 946657438, 946658337, 946659237, 946660136, 
    946661063, 946662073, 946664772, 946665682, 946666639, 946667669, 
    946668539, 946670342, 946672267, 946673160, 946678021, 946679041, 
    946684031, 946684967, 946687805, 946688547, 946688712, 946690589, 
    946691167, 946692535, 946692942, 946693258, 946694168, 946694545, 
    946696811, 946697008, 946697910, 946698667, 946698759, 946698789, 
    946699561, 946700460, 946700611, 946701079, 946701364, 946702258, 
    946702579, 946703165, 946703916, 946704055, 946704642, 946704660, 
    946705863, 946706641, 946706773, 946706992, 946707673, 946708548, 
    946709528, 946709829, 946710545, 946710546, 946710569, 946714767, 
    946716356, 946722219, 946728131, 946739875, 946740795, 946742576, 
    946749185, 946751152, 946752059, 946772296, 946773472, 946776116, 
    946776751, 946778209, 946779302, 946781974, 946782734, 946783064, 
    946783565, 946783880, 946785279, 946786233, 946786628, 946787777, 
    946788995, 946789165, 946789524, 946790012, 946791345, 946792439, 
    946792738, 946793811, 946794775, 946794838, 946796001, 946796001, 
    946798423, 946806830, 946812614, 946814489, 946820983, 946821268, 
    946823199, 946824104, 946826555, 946828880, 946830248, 946832816, 
    946839739, 946839794, 946839965, 946840682, 946840685, 946843606, 
    946844554, 946845477, 946845477, 946845639, 946849265, 946852925, 
    946853884, 946857737, 946858522, 946858633, 946859582, 946860481, 
    946861392, 946862522, 946864216, 946867763, 946868446, 946869219, 
    946870084, 946872905, 946873951, 946874497, 946874861, 946875271, 
    946876044, 946877591, 946878911, 946879707, 946880106, 946881732, 
    946882020, 946882948, 946883567, 946884924, 946887200, 946896784, 
    946898586, 946901243, 946902261, 946907060, 946909202, 946912348, 
    946913876, 946914295, 946917192, 946920238, 946926075, 946927174, 
    946943736, 946948433, 946952144, 946952518, 946953617, 946954139, 
    946954652, 946955177, 946955626, 946956623, 946957496, 946958343, 
    946958389, 946960195, 946960625, 946961260, 946961339, 946962995, 
    946964074, 946964118, 946966134, 946966502, 946966886, 946968408, 
    946970127, 946970129, 946972322, 946973321, 946974754, 946981382, 
    946987496, 946991133, 946992076, 947002878, 947033828, 947034961, 
    947037055, 947039711, 947039826, 947042697, 947043197, 947045518, 
    947045836, 947046064, 947046746, 947048020, 947048748, 947049158, 
    947051251, 947052024, 947052889, 947054754, 947055027, 947057211, 
    947058895, 947059577, 947061306, 947119101, 947125094, 947125411, 
    947125981, 947127424, 947128548, 947129850, 947130460, 947131043, 
    947131497, 947133283, 947136463, 947139449, 947139450, 947140506, 
    947141431, 947142727, 947144899, 947146595, 947150831, 947151462, 
    947152432, 947153370, 947155678, 947156575, 947162548, 947169688, 
    947170564, 947171555, 947172422, 947174355, 947175612, 947176315, 
    947177247, 947178093, 947178116, 947179271, 947180257, 947180402, 
    947180461, 947181383, 947181525, 947182474, 947182757, 947184124, 
    947186336, 947186717, 947188512, 947188811, 947190223, 947191879, 
    947192252, 947192288, 947192862, 947193784, 947194414, 947194750, 
    947194752, 947195738, 947196387, 947196713, 947197860, 947198852, 
    947200785, 947201695, 947202195, 947202686, 947205187, 947205385, 
    947211002, 947211286, 947211799, 947211989, 947213044, 947213812, 
    947215640, 947215730, 947217417, 947217810, 947218144, 947219492, 
    947221564, 947221610, 947223612, 947223809, 947224067, 947224067, 
    947225523, 947227434, 947227980, 947229754, 947230027, 947230391, 
    947231620, 947233485, 947273935, 947296921, 947300697, 947302517, 
    947303109, 947306673, 947308478, 947309843, 947310662, 947312527, 
    947315212, 947325924, 947331614, 947343867, 947344257, 947347109, 
    947353118, 947353692, 947354614, 947356514, 947359087, 947359650, 
    947360459, 947362126, 947369308, 947376843, 947379683, 947380437, 
    947382659, 947384646, 947385535, 947385673, 947386128, 947387504, 
    947388913, 947389484, 947389811, 947391708, 947391847, 947392826, 
    947394843, 947395528, 947395740, 947396870, 947398020, 947398141, 
    947398611, 947400209, 947400515, 947401437, 947410480, 947411883, 
    947415596, 947416389, 947426624, 947427840, 947435765, 947439077, 
    947441035, 947441817, 947443758, 947444679, 947444679, 947445981, 
    947445981, 947447404, 947451404, 947451404, 947453053, 947453407, 
    947464718, 947465440, 947468474, 947470432, 947471330, 947472310, 
    947474626, 947475217, 947475381, 947476746, 947477248, 947477248, 
    947481065, 947481065, 947482598, 947483023, 947483403, 947485755, 
    947487435, 947487536, 947488954, 947489356, 947493504, 947495135, 
    947498285, 947504195, 947507177, 947508240, 947509224, 947510263, 
    947512661, 947517176, 947525338, 947532247, 947545701, 947554411, 
    947554487, 947555164, 947555652, 947560521, 947561580, 947562043, 
    947563931, 947566029, 947567809, 947567999, 947570935, 947572207, 
    947572883, 947573875, 947574429, 947576716, 947579216, 947580382, 
    947583642, 947586367, 947588158, 947591281, 947600762, 947615639, 
    947617570, 947618520, 947628311, 947629199, 947630114, 947630996, 
    947631896, 947635497, 947636403, 947637378, 947639807, 947640405, 
    947644916, 947645568, 947645659, 947646296, 947646342, 947646751, 
    947647434, 947651938, 947652439, 947652484, 947653485, 947657489, 
    947658308, 947658490, 947658581, 947659491, 947661948, 947663404, 
    947665634, 947676700, 947677615, 947681774, 947687811, 947689684, 
    947689684, 947724841, 947725269, 947725587, 947726520, 947730929, 
    947731422, 947731422, 947736841, 947736916, 947737456, 947738858, 
    947750793, 947750793, 947753234, 947756487, 947762240, 947763132, 
    947771579, 947773554, 947774493, 947775786, 947776294, 947777890, 
    947780955, 947781903, 947790483, 947791375, 947792381, 947793383, 
    947794365, 947795279, 947796376, 947798220, 947799115, 947800015, 
    947807475, 947808358, 947810161, 947810244, 947811262, 947812090, 
    947812335, 947812885, 947815988, 947817054, 947817925, 947818242, 
    947821339, 947822150, 947822332, 947822762, 947823363, 947823607, 
    947823935, 947823936, 947826401, 947826504, 947827461, 947827469, 
    947827631, 947828198, 947828533, 947829477, 947829982, 947830173, 
    947830384, 947835877, 947836533, 947841933, 947846665, 947849391, 
    947852474, 947861320, 947862497, 947865788, 947867069, 947868770, 
    947871029, 947871398, 947871398, 947872066, 947873276, 947873542, 
    947874368, 947885735, 947887519, 947888400, 947896849, 947897252, 
    947901088, 947902732, 947902959, 947903824, 947906008, 947906736, 
    947906781, 947908692, 947909193, 947909739, 947912014, 947912696, 
    947912787, 947914789, 947915972, 947917337, 947918065, 947918793, 
    947920613, 947921751, 947923252, 947971793, 947982359, 947984459, 
    947985360, 947987310, 947988240, 947988528, 947989135, 947990134, 
    947991697, 947992973, 947995066, 947995596, 947996484, 947996922, 
    947997973, 947997973, 948000116, 948001434, 948002325, 948002516, 
    948002516, 948003917, 948004281, 948006061, 948007415, 948018436, 
    948021235, 948025659, 948031543, 948031769, 948032393, 948032686, 
    948033603, 948035466, 948037773, 948038845, 948041336, 948041686, 
    948044439, 948048118, 948051041, 948054296, 948060350, 948061257, 
    948070903, 948074281, 948075068, 948075304, 948076578, 948077381, 
    948080783, 948081055, 948081523, 948082855, 948083047, 948085516, 
    948086594, 948087006, 948087124, 948089480, 948091310, 948092107, 
    948092870, 948093405, 948093501, 948095192, 948097256, 948098770, 
    948110493, 948116460, 948117372, 948118329, 948121135, 948131667, 
    948132620, 948133575, 948145655, 948146686, 948149459, 948154254, 
    948156687, 948160035, 948160654, 948160985, 948161592, 948161651, 
    948162539, 948164458, 948165846, 948166775, 948167837, 948168648, 
    948169083, 948170162, 948171578, 948172373, 948172752, 948172862, 
    948173772, 948174288, 948176181, 948176278, 948177737, 948178807, 
    948178921, 948180324, 948182523, 948184956, 948186240, 948187212, 
    948208182, 948240874, 948243552, 948246610, 948252186, 948252551, 
    948256440, 948258024, 948261273, 948262306, 948264423, 948267179, 
    948267463, 948268977, 948270776, 948275476, 948278226, 948290015, 
    948291071, 948295740, 948298410, 948299573, 948313328, 948324281, 
    948326505, 948331436, 948331534, 948332455, 948332982, 948334505, 
    948337392, 948337725, 948338307, 948338406, 948339013, 948340530, 
    948340649, 948343398, 948344176, 948344612, 948346366, 948346572, 
    948347370, 948349048, 948350222, 948350627, 948352421, 948352667, 
    948356256, 948356783, 948358661, 948360329, 948375847, 948416446, 
    948417126, 948417790, 948420123, 948422438, 948423118, 948423937, 
    948423957, 948425087, 948426085, 948428538, 948429396, 948429822, 
    948429896, 948431254, 948431539, 948434454, 948434454, 948436101, 
    948436101, 948437432, 948437840, 948438656, 948439556, 948442260, 
    948443534, 948460187, 948507013, 948507599, 948509383, 948509696, 
    948509723, 948510986, 948513210, 948515218, 948515312, 948515522, 
    948515757, 948516695, 948519342, 948519600, 948521008, 948521436, 
    948521674, 948523037, 948527026, 948527504, 948527847, 948529108, 
    948531903, 948538692, 948539263, 948541742, 948550759, 948552741, 
    948556690, 948559189, 948563340, 948564842, 948564842, 948565448, 
    948566285, 948566595, 948567571, 948569159, 948588762, 948592200, 
    948592218, 948594455, 948600318, 948600350, 948600746, 948601182, 
    948604375, 948605989, 948606773, 948607411, 948607748, 948607933, 
    948609612, 948610775, 948612135, 948612199, 948613369, 948613835, 
    948614156, 948615062, 948615968, 948620154, 948625736, 948626725, 
    948629443, 948629579, 948635384, 948638518, 948641482, 948641862, 
    948642306, 948643263, 948644552, 948646037, 948647814, 948649828, 
    948651222, 948651550, 948662483, 948674483, 948677064, 948680438, 
    948681191, 948681248, 948682921, 948683355, 948684656, 948685256, 
    948686168, 948686184, 948687209, 948687435, 948689043, 948690694, 
    948691246, 948692950, 948693524, 948694964, 948695691, 948697279, 
    948698968, 948699238, 948700220, 948701122, 948704699, 948708428, 
    948709336, 948710349, 948711361, 948712271, 948717277, 948718320, 
    948719352, 948720237, 948724090, 948724283, 948725804, 948726495, 
    948730034, 948730428, 948731906, 948732501, 948738368, 948741115, 
    948744237, 948745149, 948746936, 948747875, 948752522, 948756540, 
    948757506, 948758404, 948759886, 948760321, 948761272, 948762027, 
    948763187, 948766155, 948768180, 948769064, 948769174, 948770092, 
    948770593, 948771052, 948772017, 948772534, 948772779, 948772986, 
    948774022, 948775025, 948775264, 948775973, 948776578, 948776959, 
    948777838, 948778298, 948778811, 948781014, 948781176, 948782339, 
    948784511, 948784769, 948790423, 948797982, 948804434, 948807401, 
    948808565, 948809790, 948810447, 948815974, 948816251, 948817254, 
    948829745, 948845663, 948849555, 948851729, 948855530, 948857484, 
    948857641, 948858691, 948859760, 948861475, 948863381, 948865929, 
    948866303, 948867592, 948869242, 948870593, 948871697, 948873730, 
    948875532, 948884346, 948885248, 948889015, 948895004, 948895773, 
    948931439, 948937296, 948937881, 948938203, 948938290, 948942955, 
    948943630, 948943630, 948943925, 948944361, 948944361, 948945354, 
    948946710, 948948837, 948950020, 948950049, 948950392, 948952675, 
    948952688, 948954569, 948955964, 948957672, 948958803, 948960605, 
    948962283, 948965965, 948973658, 948979438, 948993817, 948998523, 
    949011032, 949016665, 949022654, 949023119, 949023141, 949025191, 
    949026291, 949027159, 949027949, 949028855, 949029031, 949029708, 
    949032207, 949033104, 949033724, 949034798, 949034798, 949035215, 
    949036141, 949036427, 949037780, 949039702, 949040795, 949041921, 
    949042203, 949044186, 949045608, 949048010, 949051937, 949056128, 
    949057196, 949058187, 949059067, 949062784, 949064044, 949064693, 
    949066890, 949069871, 949072001, 949072969, 949082999, 949087496, 
    949095601, 949096501, 949097398, 949098300, 949102804, 949107694, 
    949108794, 949111281, 949113552, 949113552, 949114703, 949115607, 
    949117022, 949118283, 949118920, 949119425, 949119637, 949123127, 
    949124797, 949125234, 949127468, 949127637, 949129067, 949130755, 
    949131362, 949132256, 949133583, 949133607, 949137046, 949139116, 
    949140922, 949156618, 949157520, 949158430, 949194511, 949198054, 
    949198472, 949200537, 949201179, 949201179, 949202259, 949203881, 
    949204250, 949204434, 949206511, 949206884, 949207199, 949208151, 
    949209862, 949209965, 949210490, 949211335, 949212235, 949212843, 
    949212979, 949214162, 949215800, 949216104, 949218576, 949219258, 
    949220259, 949222261, 949257018, 949257897, 949258840, 949264623, 
    949266425, 949277216, 949285986, 949288625, 949289080, 949292129, 
    949293175, 949294540, 949294904, 949294950, 949297900, 949299131, 
    949299586, 949300456, 949301330, 949301397, 949304656, 949305016, 
    949305560, 949305635, 949307350, 949307386, 949309215, 949311060, 
    949311971, 949313043, 949313953, 949314984, 949316000, 949317082, 
    949318092, 949323719, 949329668, 949330145, 949344536, 949355644, 
    949356570, 949366191, 949368248, 949371933, 949374085, 949380072, 
    949380563, 949381497, 949382404, 949383497, 949384393, 949384592, 
    949384607, 949384977, 949385276, 949386383, 949390571, 949390924, 
    949393157, 949404013, 949414156, 949420059, 949422324, 949423704, 
    949426111, 949427823, 949428354, 949428357, 949429178, 949429446, 
    949430051, 949431037, 949433119, 949434071, 949434071, 949434646, 
    949435911, 949436031, 949440733, 949446728, 949447620, 949448532, 
    949451645, 949453330, 949456096, 949457473, 949458127, 949458774, 
    949459439, 949459852, 949461137, 949463719, 949463719, 949463719, 
    949464269, 949465672, 949468514, 949469668, 949469764, 949470401, 
    949471073, 949471384, 949474273, 949475349, 949475606, 949475818, 
    949476519, 949477285, 949478660, 949480748, 949489412, 949492751, 
    949494322, 949496759, 949497845, 949498490, 949501192, 949501441, 
    949502641, 949507606, 949509138, 949510975, 949511888, 949512930, 
    949513438, 949513680, 949513916, 949514194, 949514919, 949514920, 
    949517883, 949518929, 949519634, 949519967, 949520315, 949520626, 
    949521014, 949521218, 949524261, 949524601, 949525174, 949525493, 
    949526657, 949527292, 949535001, 949535943, 949537520, 949537774, 
    949538973, 949543307, 949543307, 949544053, 949548108, 949548878, 
    949549604, 949549807, 949550012, 949550752, 949553828, 949553974, 
    949554535, 949555062, 949555445, 949556259, 949556308, 949556418, 
    949558155, 949559089, 949559749, 949559773, 949562104, 949562111, 
    949562617, 949563167, 949564078, 949566000, 949567069, 949568133, 
    949568671, 949583472, 949589369, 949599318, 949610163, 949613964, 
    949614841, 949616788, 949620693, 949624161, 949628384, 949629052, 
    949629271, 949629863, 949630016, 949632775, 949634233, 949634791, 
    949634923, 949635864, 949636081, 949638560, 949639967, 949641002, 
    949641617, 949641838, 949642989, 949644430, 949644461, 949645995, 
    949646960, 949647488, 949647852, 949650582, 949652084, 949700591, 
    949704176, 949705162, 949713800, 949714619, 949719260, 949719624, 
    949720625, 949720989, 949721353, 949721711, 949722599, 949725163, 
    949725800, 949726710, 949727029, 949727438, 949729713, 949731169, 
    949731806, 949732671, 949733262, 949735719, 949737357, 949738995, 
    949847645, 949848550, 949848958, 949850292, 949851425, 949855061, 
    949856349, 949859770, 949860053, 949860146, 949861586, 949861587, 
    949863100, 949864496, 949866036, 949867596, 949869038, 949872064, 
    949872064, 949872927, 949880223, 949880533, 949881526, 949882574, 
    949883719, 949885432, 949886174, 949887283, 949889936, 949889936, 
    949889999, 949891404, 949892066, 949892066, 949892817, 949895269, 
    949895662, 949897139, 949897558, 949898108, 949898283, 949898735, 
    949899356, 949899966, 949901480, 949901509, 949903123, 949903916, 
    949904024, 949904666, 949906182, 949906629, 949907569, 949909373, 
    949910058, 949910941, 949913047, 949915919, 949916984, 949919054, 
    949921502, 949927438, 949930892, 949932020, 949933028, 949933472, 
    949933954, 949935720, 949935985, 949938893, 949939316, 949942207, 
    949942523, 949943406, 949944440, 949944984, 949945467, 949946520, 
    949946874, 949947432, 949948158, 949949158, 949950448, 949951188, 
    949951381, 949952280, 949953024, 949953351, 949954350, 949954917, 
    949955796, 949957074, 949957465, 949959128, 949962034, 949963476, 
    949965857, 949968537, 949970866, 949972085, 949972789, 949974436, 
    949977648, 949978425, 949978858, 949979356, 949980238, 949980979, 
    949983869, 949983998, 949984666, 949985565, 949986131, 949986610, 
    949988325, 949988745, 949990319, 949991041, 949992681, 949992686, 
    949992965, 949994484, 949994604, 949994820, 949996845, 949997098, 
    949998778, 949999500, 950000390, 950000416, 950000595, 950002246, 
    950003256, 950006203, 950009452, 950011602, 950012721, 950013600, 
    950017797, 950021693, 950023836, 950031149, 950032040, 950050268, 
    950055665, 950057364, 950059417, 950060074, 950061810, 950063329, 
    950064728, 950065226, 950065617, 950067412, 950069447, 950070153, 
    950070312, 950071366, 950071802, 950073190, 950073502, 950076128, 
    950076516, 950077229, 950077863, 950079316, 950079361, 950082347, 
    950082426, 950084080, 950113218, 950114097, 950115000, 950115896, 
    950140064, 950141888, 950142809, 950149015, 950150006, 950151847, 
    950155159, 950155811, 950156240, 950156968, 950157188, 950157844, 
    950158509, 950158976, 950159883, 950161660, 950162009, 950162816, 
    950163581, 950163857, 950164465, 950167436, 950168227, 950169028, 
    950169028, 950193452, 950194469, 950195391, 950196302, 950200796, 
    950202743, 950203746, 950210280, 950227254, 950228173, 950229060, 
    950229075, 950229956, 950232150, 950234698, 950235076, 950236171, 
    950238130, 950241114, 950241114, 950241844, 950242110, 950242432, 
    950243801, 950246603, 950247002, 950247509, 950248031, 950248234, 
    950249750, 950252681, 950253845, 950254066, 950254226, 950255721, 
    950259822, 950271452, 950277458, 950278777, 950314051, 950314551, 
    950320059, 950320605, 950325838, 950326566, 950326884, 950327248, 
    950327248, 950329114, 950331662, 950331935, 950332845, 950332890, 
    950333209, 950333209, 950334938, 950337895, 950338077, 950339300, 
    950339389, 950341097, 950356319, 950364285, 950370187, 950372975, 
    950373845, 950384817, 950385770, 950386743, 950387750, 950393471, 
    950395294, 950400178, 950406214, 950410825, 950411371, 950412250, 
    950412645, 950412963, 950414309, 950414309, 950417016, 950417361, 
    950418579, 950418672, 950418766, 950420054, 950422853, 950422922, 
    950423266, 950424546, 950424957, 950425680, 950426325, 950426579, 
    950427482, 950428395, 950429283, 950433058, 950433971, 950447569, 
    950451463, 950460363, 950468058, 950470886, 950479556, 950486548, 
    950486879, 950487654, 950488645, 950489558, 950489893, 950490569, 
    950491531, 950492479, 950492926, 950493729, 950495549, 950495739, 
    950497731, 950498237, 950498785, 950501812, 950501858, 950502285, 
    950503590, 950504429, 950504569, 950505302, 950507819, 950507951, 
    950508039, 950509562, 950511279, 950513645, 950515728, 950517147, 
    950517578, 950525433, 950548579, 950556181, 950565301, 950572503, 
    950574422, 950576335, 950577630, 950580311, 950580806, 950582097, 
    950583054, 950583897, 950586683, 950586711, 950587475, 950589108, 
    950589766, 950590479, 950590579, 950590629, 950591396, 950592210, 
    950592308, 950592839, 950593195, 950593592, 950594100, 950594778, 
    950596410, 950596487, 950597116, 950598493, 950598718, 950599341, 
    950600705, 950602632, 950602632, 950602839, 950604927, 950619439, 
    950620321, 950621401, 950621746, 950623282, 950627111, 950627422, 
    950627987, 950631209, 950633035, 950633718, 950633923, 950636381, 
    950638339, 950640207, 950640207, 950640207, 950642023, 950642836, 
    950644910, 950645788, 950646602, 950646635, 950650088, 950650977, 
    950651879, 950652780, 950653678, 950654584, 950655477, 950663532, 
    950665486, 950666285, 950668988, 950669381, 950670942, 950671291, 
    950675701, 950675906, 950675963, 950676348, 950677563, 950678773, 
    950680202, 950681491, 950682109, 950682914, 950683564, 950683807, 
    950684257, 950684699, 950687523, 950687846, 950688325, 950690517, 
    950700495, 950706467, 950734678, 950738514, 950739430, 950740440, 
    950747591, 950749182, 950750449, 950754870, 950755461, 950755871, 
    950756235, 950759056, 950761149, 950761513, 950761968, 950762514, 
    950765107, 950766700, 950767473, 950767564, 950768429, 950769703, 
    950770886, 950772569, 950773707, 950777165, 950778803, 950834746, 
    950835778, 950837164, 950839002, 950839920, 950840698, 950840820, 
    950841218, 950841724, 950841769, 950844330, 950846046, 950846052, 
    950846834, 950847315, 950847362, 950848217, 950848926, 950850424, 
    950851763, 950852219, 950853299, 950853535, 950853802, 950854615, 
    950856117, 950857712, 950857892, 950859712, 950862389, 950863668, 
    950864176, 950865855, 950867660, 950868648, 950869690, 950872565, 
    950890077, 950892880, 950899698, 950903771, 950918208, 950920252, 
    950920446, 950920930, 950926210, 950926286, 950929455, 950930562, 
    950931759, 950931990, 950932481, 950932853, 950933271, 950935839, 
    950936383, 950937026, 950938224, 950939244, 950939836, 950941314, 
    950941533, 950942306, 950942907, 950945235, 950945410, 950946052, 
    950950863, 950951763, 950955358, 950958065, 950962122, 950968501, 
    950994719, 950995619, 950997417, 951004916, 951006155, 951010741, 
    951011333, 951012044, 951012549, 951012967, 951013167, 951013973, 
    951014821, 951014983, 951016396, 951016754, 951017218, 951018233, 
    951018892, 951019967, 951020497, 951021071, 951022311, 951023088, 
    951024980, 951025108, 951026853, 951026898, 951028317, 951028520, 
    951030193, 951031204, 951031216, 951032794, 951032794, 951038782, 
    951039789, 951044653, 951046181, 951047143, 951048139, 951049152, 
    951050101, 951050226, 951051002, 951056168, 951064651, 951070377, 
    951071327, 951072422, 951073471, 951080101, 951081037, 951082168, 
    951085978, 951091904, 951096035, 951097986, 951098783, 951101626, 
    951101927, 951103501, 951103974, 951104401, 951105299, 951105502, 
    951105828, 951107374, 951108019, 951109234, 951110212, 951110301, 
    951110517, 951111246, 951111456, 951111726, 951112138, 951113104, 
    951113374, 951116749, 951116757, 951118007, 951119649, 951122098, 
    951122871, 951123872, 951125647, 951128464, 951129360, 951177596, 
    951180994, 951183591, 951186854, 951186854, 951189940, 951189940, 
    951190332, 951191046, 951192483, 951193094, 951193468, 951194429, 
    951195684, 951196077, 951196359, 951197071, 951198425, 951199210, 
    951201441, 951201930, 951202619, 951203029, 951204738, 951207779, 
    951208552, 951210789, 951219666, 951240383, 951264587, 951265236, 
    951265935, 951266140, 951267017, 951267984, 951269072, 951269611, 
    951272039, 951272039, 951275268, 951276141, 951276162, 951277598, 
    951278039, 951280521, 951280526, 951281560, 951282227, 951282227, 
    951283480, 951283662, 951286492, 951287000, 951287913, 951288238, 
    951288896, 951294151, 951294151, 951295931, 951298350, 951304285, 
    951306409, 951307461, 951320103, 951321032, 951336728, 951337685, 
    951341370, 951354973, 951355381, 951355670, 951355858, 951356557, 
    951357996, 951359049, 951360234, 951360969, 951362009, 951362705, 
    951362984, 951363328, 951365010, 951366099, 951367143, 951367372, 
    951367631, 951368699, 951368822, 951372045, 951373137, 951373696, 
    951374924, 951377123, 951377740, 951378121, 951379115, 951379208, 
    951381100, 951388782, 951400294, 951401276, 951405421, 951406306, 
    951406315, 951408403, 951411394, 951412193, 951412194, 951423201, 
    951424667, 951430136, 951434783, 951440764, 951441707, 951441755, 
    951442085, 951446631, 951447359, 951449679, 951452910, 951453319, 
    951453638, 951453865, 951455731, 951456823, 951459143, 951459553, 
    951459735, 951461646, 951463011, 951464467, 951465650, 951466241, 
    951508041, 951508923, 951509821, 951510719, 951511655, 951521350, 
    951526615, 951526748, 951527320, 951528710, 951530654, 951532454, 
    951532454, 951532458, 951536434, 951538493, 951539020, 951539020, 
    951539559, 951540059, 951540466, 951542032, 951543064, 951544516, 
    951544922, 951545004, 951545229, 951545826, 951546304, 951548088, 
    951548595, 951551250, 951551338, 951551364, 951552077, 951552254, 
    951553135, 951558556, 951559455, 951560350, 951561251, 951562190, 
    951563202, 951565601, 951569606, 951576916, 951577827, 951579658, 
    951581475, 951582477, 951583488, 951585444, 951586498, 951587599, 
    951592566, 951594773, 951595679, 951596783, 951598696, 951601665, 
    951611512, 951612383, 951615423, 951616322, 951617971, 951618116, 
    951618900, 951619022, 951623168, 951624140, 951624695, 951627453, 
    951629346, 951630385, 951630843, 951630843, 951633395, 951636120, 
    951636740, 951659950, 951662477, 951662810, 951666191, 951666863, 
    951667961, 951697905, 951697905, 951698469, 951703870, 951704006, 
    951706786, 951708074, 951708595, 951709299, 951709477, 951709999, 
    951710445, 951713833, 951713933, 951715316, 951715453, 951716453, 
    951718413, 951719401, 951719759, 951721288, 951721400, 951722655, 
    951723006, 951725726, 951725929, 951727671, 951739271, 951743819, 
    951757806, 951759612, 951761408, 951762295, 951763213, 951766796, 
    951767696, 951769501, 951771297, 951772196, 951783060, 951786674, 
    951789413, 951789554, 951790389, 951792192, 951793052, 951793899, 
    951795715, 951796443, 951797937, 951799318, 951799318, 951799566, 
    951800767, 951802151, 951803516, 951804976, 951805214, 951805682, 
    951807115, 951808016, 951809580, 951812789, 951820746, 951823316, 
    951836914, 951841718, 951842774, 951843844, 951869261, 951870107, 
    951872127, 951872438, 951875349, 951875974, 951877880, 951878267, 
    951878318, 951878439, 951880068, 951881479, 951881800, 951881941, 
    951882843, 951884033, 951884103, 951884182, 951885540, 951885755, 
    951886451, 951887350, 951887416, 951887993, 951888653, 951890048, 
    951890126, 951890126, 951891734, 951892022, 951893719, 951893835, 
    951895619, 951896184, 951898019, 951898316, 951899216, 951900114, 
    951915607, 951955196, 951960974, 951962749, 951962931, 951966844, 
    951968573, 951968800, 951969255, 951971030, 951973214, 951973487, 
    951974852, 951974897, 951975261, 952016087, 952017302, 952017844, 
    952018455, 952018972, 952020700, 952021737, 952023353, 952023457, 
    952023663, 952024524, 952025159, 952026660, 952029921, 952030264, 
    952031057, 952032531, 952033393, 952034350, 952034957, 952035240, 
    952035516, 952035516, 952036145, 952036191, 952036799, 952038578, 
    952039242, 952040719, 952041258, 952041608, 952042880, 952044690, 
    952046598, 952047561, 952047904, 952048723, 952050486, 952052819, 
    952053225, 952053226, 952053651, 952054889, 952056512, 952058964, 
    952059015, 952059283, 952059802, 952060612, 952062292, 952065303, 
    952065303, 952066557, 952068342, 952071257, 952071591, 952074225, 
    952074487, 952082007, 952088739, 952094415, 952096522, 952100740, 
    952103409, 952103940, 952105730, 952106647, 952107552, 952108728, 
    952109310, 952109310, 952109952, 952111598, 952132394, 952132969, 
    952133223, 952134027, 952135661, 952137693, 952138466, 952138467, 
    952139044, 952139599, 952141588, 952143915, 952144277, 952144607, 
    952144845, 952144845, 952145515, 952147233, 952150062, 952150223, 
    952153612, 952155765, 952156275, 952157059, 952166969, 952178957, 
    952181186, 952191848, 952195951, 952214817, 952218380, 952218968, 
    952223362, 952228036, 952228482, 952229036, 952229644, 952230004, 
    952230307, 952230533, 952230673, 952230903, 952232424, 952234377, 
    952235602, 952236540, 952236540, 952238648, 952240168, 952242654, 
    952243122, 952251668, 952253466, 952254376, 952268378, 952280686, 
    952302566, 952303887, 952305578, 952306585, 952307458, 952308381, 
    952308428, 952309687, 952310159, 952312938, 952314119, 952314351, 
    952316086, 952316112, 952316275, 952317616, 952319780, 952320696, 
    952320696, 952321896, 952322371, 952323396, 952326810, 952329750, 
    952478465, 952481345, 952481923, 952484221, 952486226, 952487371, 
    952487699, 952487968, 952490224, 952492438, 952493433, 952493696, 
    952493720, 952494057, 952496337, 952496754, 952498765, 952500006, 
    952500006, 952500382, 952504450, 952505857, 952506286, 952512453, 
    952513322, 952514273, 952516197, 952517471, 952523115, 952525231, 
    952529255, 952531052, 952533789, 952538513, 952539561, 952541425, 
    952545665, 952561346, 952561539, 952561809, 952563208, 952566860, 
    952569075, 952571425, 952572315, 952572954, 952573325, 952573325, 
    952574555, 952575229, 952577495, 952578802, 952579031, 952579249, 
    952579691, 952580962, 952581878, 952583409, 952583631, 952584655, 
    952585137, 952585282, 952588226, 952589446, 952590069, 952591279, 
    952591537, 952598159, 952599063, 952609920, 952623861, 952626771, 
    952631732, 952632595, 952634398, 952635319, 952636307, 952637219, 
    952638198, 952639136, 952646649, 952646840, 952650032, 952652054, 
    952652550, 952653035, 952653923, 952656661, 952656881, 952656898, 
    952657593, 952658269, 952658687, 952659005, 952660115, 952661555, 
    952662781, 952662980, 952664085, 952664828, 952665009, 952666303, 
    952666976, 952668508, 952669021, 952670178, 952671069, 952673181, 
    952674529, 952674893, 952676375, 952682446, 952710296, 952713985, 
    952723881, 952733218, 952733939, 952738312, 952738502, 952739221, 
    952743759, 952744341, 952744751, 952744823, 952747641, 952747700, 
    952749811, 952750454, 952750763, 952751149, 952752459, 952753542, 
    952753683, 952755917, 952757002, 952757037, 952758708, 952759526, 
    952759820, 952761472, 952773902, 952774798, 952780569, 952790118, 
    952811319, 952813141, 952821415, 952822368, 952823930, 952827176, 
    952830070, 952830101, 952830548, 952832450, 952834852, 952835903, 
    952835904, 952836175, 952836470, 952836775, 952837680, 952838110, 
    952838888, 952840431, 952840432, 952841364, 952841863, 952842694, 
    952843443, 952844035, 952844141, 952844936, 952844939, 952846395, 
    952848488, 952849398, 952850945, 953036041, 953036511, 953037030, 
    953042335, 953043445, 953044428, 953045311, 953048108, 953049087, 
    953054060, 953054953, 953054957, 953055837, 953057086, 953057291, 
    953058145, 953058897, 953059128, 953059806, 953060747, 953060805, 
    953060977, 953061747, 953062653, 953063369, 953063550, 953063754, 
    953064416, 953064750, 953065328, 953066270, 953066403, 953069666, 
    953070341, 953070993, 953072721, 953072854, 953073749, 953074638, 
    953075264, 953085680, 953086627, 953086957, 953088586, 953090220, 
    953090336, 953091690, 953093063, 953093609, 953093837, 953094701, 
    953094730, 953095626, 953096588, 953096628, 953097688, 953098527, 
    953098878, 953099533, 953100268, 953102024, 953103196, 953105155, 
    953106644, 953109363, 953113320, 953114225, 953115307, 953120925, 
    953128796, 953129703, 953131197, 953131885, 953135122, 953137162, 
    953138968, 953139026, 953139950, 953140018, 953142012, 953143092, 
    953144257, 953146290, 953148733, 953149681, 953150064, 953151781, 
    953154723, 953155671, 953156270, 953157611, 953157914, 953164081, 
    953165215, 953166209, 953167214, 953167215, 953167700, 953168270, 
    953169412, 953175701, 953176182, 953176221, 953178724, 953180530, 
    953181450, 953181477, 953181480, 953182100, 953185239, 953185642, 
    953187512, 953187537, 953188392, 953190223, 953191205, 953193095, 
    953193784, 953193988, 953196079, 953205124, 953207171, 953208155, 
    953211506, 953213996, 953214898, 953216988, 953217299, 953222934, 
    953223383, 953224841, 953232953, 953240410, 953249089, 953250005, 
    953251006, 953252150, 953252462, 953256863, 953258478, 953258900, 
    953260713, 953264171, 953265955, 953266302, 953266624, 953266624, 
    953269411, 953271332, 953272325, 953272501, 953272709, 953276714, 
    953276789, 953277373, 953277834, 953278493, 953280173, 953282945, 
    953283211, 953287932, 953294847, 953302152, 953302523, 953307651, 
    953308636, 953313116, 953313929, 953314564, 953314678, 953315018, 
    953315653, 953315804, 953317623, 953320280, 953320719, 953324166, 
    953332530, 953333401, 953335267, 953336181, 953338348, 953341565, 
    953344271, 953349983, 953350200, 953350938, 953351369, 953354714, 
    953356654, 953357566, 953357566, 953361889, 953362926, 953363790, 
    953369529, 953386228, 953388145, 953390089, 953392534, 953394016, 
    953394802, 953398354, 953399554, 953400168, 953400478, 953405697, 
    953406110, 953406474, 953406731, 953406989, 953430002, 953430103, 
    953430555, 953435169, 953436598, 953441264, 953441783, 953442085, 
    953442235, 953442584, 953445494, 953446657, 953447275, 953448088, 
    953448422, 953448455, 953451596, 953453141, 953454751, 953462078, 
    953463002, 953464098, 953466973, 953470958, 953473047, 953475090, 
    953476999, 953480183, 953483241, 953485931, 953486288, 953486288, 
    953492367, 953492502, 953494307, 953495215, 953496238, 953497198, 
    953497484, 953497912, 953498095, 953498167, 953498167, 953514991, 
    953515674, 953520178, 953520269, 953520952, 953521543, 953521862, 
    953522104, 953526093, 953526139, 953526139, 953526912, 953527686, 
    953527777, 953528050, 953530666, 953531872, 953532509, 953533009, 
    953533737, 953533919, 953536513, 953538242, 953540001, 953540517, 
    953624962, 953625951, 953644499, 953651403, 953651749, 953655538, 
    953657250, 953658095, 953659622, 953661318, 953661345, 953662500, 
    953663216, 953663771, 953665883, 953667313, 953667352, 953669942, 
    953671471, 953673506, 953674914, 953676226, 953678909, 953681187, 
    953682672, 953686508, 953686945, 953689813, 953690796, 953690822, 
    953691613, 953692495, 953692499, 953692935, 953695253, 953696586, 
    953696614, 953698161, 953699223, 953699379, 953700752, 953702473, 
    953702777, 953704122, 953705263, 953707303, 953708849, 953710315, 
    953711400, 953713050, 953714739, 953716457, 953716692, 953718488, 
    953719383, 953724880, 953724907, 953744036, 953748697, 953749615, 
    953751649, 953752807, 953754724, 953755736, 953757539, 953760307, 
    953762491, 953764610, 953765561, 953772637, 953773031, 953773436, 
    953777887, 953778540, 953779232, 953779812, 953781474, 953781858, 
    953783332, 953784775, 953784995, 953786025, 953786049, 953787160, 
    953787262, 953787426, 953788080, 953788985, 953789261, 953790786, 
    953791169, 953791720, 953791942, 953792252, 953792651, 953793505, 
    953793644, 953795590, 953797159, 953799382, 953800311, 953801468, 
    953815280, 953821005, 953835240, 953842228, 953843129, 953846935, 
    953858757, 953864390, 953864390, 953864932, 953866272, 953868722, 
    953870385, 953870664, 953870691, 953871668, 953872614, 953872802, 
    953873141, 953874396, 953876358, 953876678, 953877274, 953878462, 
    953878601, 953878755, 953880615, 953882231, 953883169, 953883267, 
    953891996, 953893942, 953899953, 953905843, 953908305, 953911674, 
    953914289, 953916351, 953917708, 953920298, 953920747, 953921876, 
    953944079, 953945399, 953948857, 953950085, 953950631, 953951223, 
    953952133, 953953680, 953954924, 953956046, 953956501, 953957472, 
    953957911, 953959549, 953961051, 953962416, 953962461, 953963144, 
    953963872, 953965328, 954043199, 954044825, 954045571, 954048270, 
    954048270, 954049163, 954050538, 954051209, 954051488, 954054133, 
    954055423, 954056609, 954057037, 954057387, 954057483, 954058375, 
    954059304, 954060192, 954060454, 954061996, 954062891, 954063264, 
    954067109, 954070205, 954074924, 954077888, 954078801, 954079669, 
    954080678, 954080823, 954081855, 954082748, 954083652, 954084769, 
    954085716, 954085717, 954085843, 954086575, 954086674, 954087640, 
    954088575, 954091257, 954091806, 954091964, 954092159, 954092771, 
    954092892, 954093961, 954094315, 954098057, 954098263, 954098291, 
    954099365, 954100441, 954106361, 954107511, 954115916, 954117426, 
    954118364, 954119601, 954120476, 954121221, 954121627, 954123488, 
    954127459, 954127459, 954129580, 954130003, 954130363, 954130613, 
    954133321, 954133921, 954134305, 954135825, 954136280, 954138690, 
    954140251, 954140559, 954142050, 954142050, 954142982, 954143891, 
    954146226, 954153692, 954160236, 954161104, 954170653, 954171217, 
    954171862, 954177885, 954177909, 954182537, 954183895, 954184057, 
    954184219, 954185993, 954186609, 954187679, 954188845, 954188845, 
    954190165, 954190283, 954206416, 954207262, 954207801, 954207892, 
    954208537, 954212411, 954213107, 954213851, 954213851, 954214518, 
    954218094, 954218233, 954219576, 954219613, 954219640, 954220548, 
    954221107, 954224131, 954224154, 954225485, 954225822, 954226515, 
    954228501, 954230554, 954231516, 954231976, 954242157, 954243958, 
    954243979, 954249582, 954251153, 954255896, 954257050, 954258300, 
    954261581, 954261740, 954262172, 954263181, 954267770, 954273197, 
    954274259, 954292835, 954292835, 954293687, 954297099, 954298816, 
    954299122, 954299254, 954299520, 954300330, 954303029, 954304918, 
    954304918, 954305297, 954305516, 954306323, 954310482, 954311222, 
    954311222, 954312768, 954314655, 954318386, 954318797, 954328634, 
    954334475, 954334607, 954335566, 954337611, 954340205, 954341376, 
    954342992, 954343200, 954344105, 954346353, 954346474, 954348870, 
    954350408, 954354336, 954355096, 954355097, 954356024, 954362629, 
    954364550, 954369579, 954375365, 954376258, 954377173, 954378745, 
    954379149, 954382000, 954382027, 954383731, 954383784, 954384525, 
    954385151, 954385725, 954387935, 954389532, 954389986, 954391017, 
    954391079, 954391490, 954393842, 954395731, 954395783, 954397298, 
    954397651, 954398330, 954400475, 954401915, 954403704, 954413102, 
    954416212, 954419106, 954424696, 954427296, 954428618, 954430670, 
    954431595, 954434535, 954434875, 954436764, 954437643, 954438655, 
    954441377, 954449706, 954450596, 954453381, 954457982, 954458905, 
    954464407, 954466773, 954468184, 954469048, 954470140, 954470641, 
    954470732, 954472597, 954474144, 954474827, 954476328, 954476556, 
    954476783, 954478376, 954479741, 954480378, 954480833, 954482516, 
    954482653, 954485519, 954486930, 954488477, 954488750, 954567725, 
    954568480, 954569460, 954570374, 954570421, 954570506, 954572011, 
    954572235, 954573626, 954574768, 954576633, 954578276, 954579961, 
    954580170, 954585000, 954585911, 954588259, 954593972, 954595806, 
    954598851, 954599980, 954600128, 954605516, 954605913, 954605954, 
    954606418, 954607164, 954609813, 954611384, 954612095, 954612401, 
    954613174, 954616002, 954617280, 954618023, 954618710, 954619018, 
    954620246, 954621813, 954635743, 954636642, 954641662, 954642361, 
    954643178, 954643832, 954645470, 954646932, 954648116, 954648116, 
    954648383, 954649246, 954649698, 954650173, 954651075, 954652901, 
    954654140, 954654272, 954655053, 954657238, 954658722, 954660344, 
    954661257, 954661798, 954663467, 954665156, 954671522, 954672500, 
    954672765, 954673408, 954674281, 954679910, 954685239, 954696121, 
    954700680, 954702874, 954703741, 954720520, 954721404, 954721543, 
    954722173, 954723122, 954727095, 954727407, 954727596, 954727735, 
    954730660, 954732104, 954733189, 954733836, 954733836, 954733953, 
    954736313, 954738111, 954738938, 954739456, 954739819, 954739819, 
    954739891, 954740786, 954740855, 954741665, 954742650, 954742674, 
    954744548, 954745980, 954746921, 954748490, 954750109, 954752033, 
    954754266, 954758140, 954759058, 954759977, 954761016, 954761961, 
    954762961, 954763885, 954771624, 954772560, 954773634, 954774616, 
    954775049, 954776855, 954777473, 954780088, 954807306, 954812220, 
    954813084, 954818271, 954818317, 954819090, 954905065, 954905286, 
    954907049, 954908305, 954908794, 954909333, 954911528, 954912875, 
    954914419, 954914838, 954916800, 954918710, 954920546, 954920654, 
    954932355, 954937806, 954938081, 954938835, 954943728, 954948691, 
    954950013, 954952590, 954955244, 954956300, 954958766, 954960880, 
    954961509, 954962341, 954962478, 954964148, 954964366, 954964780, 
    954967229, 954967427, 954968677, 954970298, 954982458, 954984542, 
    954987288, 954987970, 954990788, 954990900, 954992317, 954993327, 
    954993491, 954993895, 954996394, 954996573, 954997008, 954997878, 
    954999395, 954999401, 955000256, 955002400, 955002797, 955003923, 
    955005241, 955005567, 955009237, 955010304, 955010351, 955011196, 
    955011739, 955014843, 955026284, 955040610, 955042520, 955048379, 
    955051202, 955058658, 955067201, 955067201, 955070240, 955070650, 
    955070967, 955071398, 955072932, 955076102, 955077336, 955077933, 
    955078904, 955078904, 955082434, 955082935, 955084076, 955084733, 
    955084733, 955087852, 955088721, 955088812, 955090838, 955094665, 
    955095206, 955112937, 955119120, 955120141, 955122309, 955125138, 
    955126085, 955126626, 955128321, 955128348, 955152118, 955156395, 
    955156681, 955157579, 955158069, 955158346, 955162116, 955162300, 
    955162452, 955164089, 955168185, 955168211, 955168211, 955168211, 
    955170112, 955170196, 955172663, 955174186, 955174209, 955175766, 
    955176005, 955178862, 955180018, 955180294, 955182149, 955197495, 
    955203492, 955206021, 955207089, 955215838, 955230395, 955241475, 
    955241860, 955244752, 955245661, 955246558, 955246878, 955247469, 
    955247584, 955248431, 955248717, 955252883, 955253599, 955253756, 
    955253982, 955254851, 955254905, 955257641, 955258139, 955259132, 
    955259132, 955259707, 955260042, 955261207, 955264311, 955265388, 
    955267230, 955272297, 955273124, 955282224, 955288048, 955291961, 
    955423997, 955424562, 955425343, 955425476, 955425476, 955426742, 
    955427672, 955427899, 955429658, 955430759, 955431450, 955431450, 
    955433645, 955433825, 955434309, 955435553, 955439751, 955443599, 
    955452357, 955453259, 955455076, 955455957, 955456900, 955457226, 
    955459004, 955460910, 955463045, 955463179, 955467889, 955469173, 
    955469235, 955482620, 955489946, 955490820, 955498806, 955498860, 
    955499297, 955500839, 955501750, 955503181, 955503533, 955504674, 
    955504817, 955506576, 955509415, 955510729, 955511560, 955512452, 
    955513694, 955515738, 955516818, 955517548, 955518367, 955519321, 
    955519321, 955520837, 955521823, 955522526, 955522742, 955523472, 
    955524373, 955527205, 955528633, 955530227, 955539312, 955541101, 
    955541686, 955542906, 955551124, 955558321, 955559271, 955560206, 
    955561085, 955584481, 955585118, 955588360, 955590418, 955591079, 
    955594354, 955594354, 955595856, 955596540, 955596973, 955597072, 
    955597239, 955599179, 955600198, 955600412, 955602709, 955602709, 
    955604817, 955606002, 955607963, 955609266, 955609267, 955611852, 
    955613946, 955614827, 955618951, 955619817, 955620717, 955622546, 
    955632058, 955634427, 955635182, 955638143, 955640761, 955640987, 
    955643731, 955647987, 955652566, 955662349, 955668204, 955670399, 
    955670930, 955671153, 955672021, 955673331, 955675937, 955676272, 
    955676936, 955680727, 955681143, 955681382, 955682498, 955682620, 
    955682621, 955684682, 955685136, 955685136, 955686684, 955686786, 
    955687539, 955688455, 955688455, 955689600, 955691215, 955691299, 
    955692632, 955694687, 955695677, 955696863, 955697118, 955698631, 
    955700736, 955712804, 955716620, 955722661, 955726165, 955728758, 
    955732353, 955772000, 955772115, 955774174, 955774290, 955775591, 
    955775848, 955776347, 955778035, 955778035, 955780365, 955781287, 
    955782390, 955782443, 955784322, 955786740, 955789861, 955790174, 
    955792935, 955793920, 955795626, 955795754, 955796689, 955801236, 
    955807191, 955811766, 955813048, 955829309, 955833930, 955843983, 
    955844885, 955847485, 955847601, 955848485, 955849173, 955850639, 
    955853823, 955853917, 955855694, 955856519, 955859855, 955859883, 
    955860993, 955861081, 955861392, 955862500, 955863110, 955865870, 
    955865957, 955867063, 955867445, 955867717, 955868463, 955869187, 
    955872250, 955873706, 955874272, 955875557, 955880008, 955891801, 
    955897507, 955897646, 955902009, 955903870, 955904607, 955905067, 
    955906960, 955909570, 955924899, 955925880, 955930557, 955933475, 
    955934124, 955934971, 955940190, 955942250, 955946118, 955946685, 
    955947296, 955948162, 955951151, 955951379, 955952067, 955952303, 
    955952778, 955954488, 955957137, 955957918, 955958702, 955970504, 
    955976240, 955976241, 955977172, 955978076, 955978976, 955982206, 
    955983343, 955988371, 955989395, 955989410, 956018999, 956042174, 
    956043307, 956043697, 956045697, 956054649, 956061117, 956066813, 
    956067964, 956068735, 956068859, 956070669, 956071565, 956072951, 
    956073361, 956074046, 956074289, 956074836, 956075359, 956078908, 
    956080327, 956080858, 956092098, 956094180, 956097191, 956099959, 
    956100836, 956101741, 956103596, 956103848, 956104872, 956105531, 
    956106454, 956110800, 956111127, 956112741, 956115596, 956116111, 
    956116664, 956117045, 956117073, 956118554, 956121567, 956122426, 
    956123453, 956124616, 956128082, 956129097, 956129260, 956130763, 
    956133888, 956135225, 956139886, 956145658, 956151581, 956179393, 
    956180279, 956183236, 956187357, 956190600, 956190661, 956196485, 
    956200519, 956200648, 956202402, 956203567, 956203778, 956206270, 
    956206643, 956206643, 956207191, 956207940, 956208515, 956209699, 
    956214733, 956215657, 956217957, 956218517, 956219877, 956221858, 
    956227800, 956229642, 956230607, 956231622, 956233676, 956235961, 
    956239407, 956240281, 956240333, 956241677, 956243877, 956244305, 
    956246580, 956250175, 956251767, 956281930, 956381876, 956382379, 
    956382897, 956384348, 956386248, 956386249, 956387799, 956388958, 
    956390422, 956392258, 956392258, 956396952, 956397996, 956398895, 
    956399817, 956400772, 956402768, 956411077, 956411378, 956417324, 
    956417689, 956419884, 956421953, 956423071, 956423694, 956424079, 
    956425802, 956427929, 956429677, 956429715, 956445062, 956449297, 
    956453330, 956453540, 956455338, 956455391, 956457936, 956459358, 
    956459358, 956459744, 956460135, 956460993, 956463602, 956465167, 
    956465764, 956465764, 956466356, 956467371, 956469568, 956471225, 
    956471774, 956473383, 956474140, 956475618, 956477458, 956477507, 
    956478021, 956479329, 956480217, 956491602, 956497329, 956498174, 
    956501409, 956503644, 956507375, 956539265, 956553259, 956554710, 
    956556395, 956556742, 956556900, 956557512, 956561051, 956562554, 
    956565790, 956568494, 956570578, 956580189, 956581405, 956585859, 
    956587405, 956588296, 956588963, 956589186, 956589607, 956591896, 
    956592097, 956595037, 956597344, 956624970, 956625035, 956628032, 
    956631241, 956631241, 956633859, 956635285, 956635895, 956637030, 
    956637106, 956637106, 956638767, 956640286, 956641201, 956643195, 
    956646113, 956647201, 956647848, 956649204, 956652171, 956653039, 
    956664681, 956670511, 956676411, 956785082, 956790409, 956794868, 
    956796233, 956801010, 956802284, 956804377, 956804650, 956806834, 
    956808518, 956808563, 956810383, 956810520, 956811930, 956812886, 
    956814433, 956814615, 956814842, 956816194, 956817699, 956820933, 
    956820992, 956822608, 956824162 ;

 z = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0 ;
}
