netcdf ATN_Trajectory {
dimensions:
	obs = < dim1 > ;
variables:
	int crs ;
		crs:epsg_code = "EPSG:4326" ;
		crs:grid_mapping_name = "latitude_longitude" ;
		crs:inverse_flattening = 298.257223563 ;
		crs:ioos_category = "Other" ;
		crs:long_name = "http://www.opengis.net/def/crs/EPSG/0/4326" ;
		crs:semi_major_axis = 6378137. ;
	double ellipse_orientation(obs) ;
		ellipse_orientation:_FillValue = -9999.9 ;
		ellipse_orientation:coordinates = "time z lon lat" ;
		ellipse_orientation:long_name = "Platform identifier" ;
		ellipse_orientation:units = "degrees" ;
		ellipse_orientation:comment = "The angle in degrees of the ellipse from true north, proceeding clockwise (0 to 360). A blank field represents 0 degrees." ;
		ellipse_orientation:instrument = "instrument_location" ;
		ellipse_orientation:platform = "platform" ;
	double error_radius(obs) ;
		error_radius:_FillValue = -9999.9 ;
		error_radius:coordinates = "time z lon lat" ;
		error_radius:long_name = "Error radius" ;
		error_radius:units = "m" ;
		error_radius:comment = "If the position is best represented as a circle, this field gives the radius of that circle in meters." ;
		error_radius:instrument = "instrument_location" ;
		error_radius:platform = "platform" ;
	string instrument_location ;
		instrument_location:long_name = "Wildlife Computers Splash 10" ;
		instrument_location:location_type = "argos / modeled" ;
		instrument_location:comment = "Location" ;
		instrument_location:manufacturer = "Wildlife Computers" ;
		instrument_location:make_model = "Splash 10" ;
		instrument_location:calibration_date = "" ;
		instrument_location:serial_number = "18A0360" ;
	string instrument_pressure ;
		instrument_pressure:long_name = "some pressure sensor" ;
		instrument_pressure:comment = "hypothetical WC pressure sensos" ;
		instrument_pressure:manufacturer = "Wildlife Computers" ;
		instrument_pressure:make_model = "WC pressure sensor" ;
		instrument_pressure:calibration_date = "" ;
		instrument_pressure:serial_number = "XXX55544XO" ;
	string instrument_tag ;
		instrument_tag:long_name = "instrument" ;
		instrument_tag:comment = "Test comment" ;
		instrument_tag:manufacturer = "Wildlife Computers" ;
		instrument_tag:make_model = "Splash 10" ;
		instrument_tag:calibration_date = "" ;
		instrument_tag:serial_number = "18A0360" ;
	double lat(obs) ;
		lat:_FillValue = -9999.9 ;
		lat:axis = "Y" ;
		lat:_CoordinateAxisType = "Lat" ;
		lat:ioos_category = "Location" ;
		lat:long_name = "Profile Location" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:valid_max = 90. ;
		lat:valid_min = -90. ;
		lat:actual_min = 50.6209 ;
		lat:actual_max = 66.8307 ;
		lat:instrument = "instrument_location" ;
		lat:platform = "platform" ;
	string location_class(obs) ;
		location_class:coordinates = "time z lon lat" ;
		location_class:long_name = "Location Quality Code" ;
		location_class:standard_name = "quality_code" ;
		location_class:ioos_category = "Quality" ;
		location_class:comment = "Quality codes from the ARGOS satellite (in meters): G,3,2,1,0,A,B,Z. See http://www.argos-system.org/manual/3-location/34_location_classes.htm" ;
		location_class:instrument = "instrument_location" ;
		location_class:platform = "platform" ;
	double lon(obs) ;
		lon:_FillValue = -9999.9 ;
		lon:axis = "X" ;
		lon:_CoordinateAxisType = "Lon" ;
		lon:ioos_category = "Location" ;
		lon:long_name = "Profile Location" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:valid_max = 180. ;
		lon:valid_min = -180. ;
		lon:actual_min = -154.258 ;
		lon:actual_max = 160.9647 ;
		lon:instrument = "instrument_location" ;
		lon:platform = "platform" ;
	double offset(obs) ;
		offset:_FillValue = -9999.9 ;
		offset:coordinates = "time z lon lat" ;
		offset:long_name = "Offset" ;
		offset:units = "m" ;
		offset:comment = "This field is non-zero if the circle or ellipse are not centered on the (Latitude, Longitude) values on this row. \"Offset\" gives the distance in meters from (Latitude, Longitude) to the center of the ellipse." ;
	double offset_orientation(obs) ;
		offset_orientation:_FillValue = -9999.9 ;
		offset_orientation:coordinates = "time z lon lat" ;
		offset_orientation:long_name = "Offset orientation" ;
		offset_orientation:units = "degrees" ;
		offset_orientation:comment = "If the \"Offset\" field is non-zero, this field is the angle in degrees from (Latitude, Longitude) to the center of the ellipse. Zero degrees is true north; a blank field represents 0 degrees." ;
	string platform ;
		platform:cf_role = "5deb0b1d6321be14905284b8" ;
		platform:long_name = "SSL2019788KOD" ;
		platform:platform_type = "animal" ;
		platform:platform_vocabulary = "https://mmisw.org/ont/ioos/platform" ;
		platform:valid_name = "Eumetopias jubatus" ;
		platform:AphiaID = 254999LL ;
		platform:scientificname = "Eumetopias jubatus" ;
		platform:authority = "(Schreber, 1776)" ;
		platform:kingdom = "Animalia" ;
		platform:phylum = "Chordata" ;
		platform:class = "Mammalia" ;
		platform:order = "Carnivora" ;
		platform:family = "Otariidae" ;
		platform:genus = "Eumetopias" ;
		platform:taxonRankID = 220LL ;
		platform:rank = "Species" ;
		platform:superdomain = "Biota" ;
		platform:subphylum = "Vertebrata" ;
		platform:superclass = "Tetrapoda" ;
		platform:subclass = "Theria" ;
		platform:suborder = "Caniformia" ;
		platform:infraorder = "Pinnipedia" ;
		platform:species = "Eumetopias jubatus" ;
	string qartod_location_flag ;
		string qartod_location_flag:_FillValue = "0" ;
		qartod_location_flag:flag_meanings = "PASS NOT_EVALUATED SUSPECT FAIL MISSING" ;
		qartod_location_flag:flag_values = "1, 2, 3, 4, 9" ;
		qartod_location_flag:ioos_category = "Other" ;
		qartod_location_flag:long_name = "" ;
		qartod_location_flag:standard_name = "" ;
	string qartod_rollup_flag2 ;
		string qartod_rollup_flag2:_FillValue = "0" ;
		qartod_rollup_flag2:flag_meanings = "PASS NOT_EVALUATED SUSPECT FAIL MISSING" ;
		qartod_rollup_flag2:flag_values = "1, 2, 3, 4, 9" ;
		qartod_rollup_flag2:ioos_category = "Other" ;
		qartod_rollup_flag2:long_name = "" ;
		qartod_rollup_flag2:standard_name = "" ;
	string qartod_speed_flag ;
		string qartod_speed_flag:_FillValue = "0" ;
		qartod_speed_flag:flag_meanings = "PASS NOT_EVALUATED SUSPECT FAIL MISSING" ;
		qartod_speed_flag:flag_values = "1, 2, 3, 4, 9" ;
		qartod_speed_flag:ioos_category = "Other" ;
		qartod_speed_flag:long_name = "" ;
		qartod_speed_flag:standard_name = "" ;
	string qartod_time_flag ;
		string qartod_time_flag:_FillValue = "0" ;
		qartod_time_flag:flag_meanings = "PASS NOT_EVALUATED SUSPECT FAIL MISSING" ;
		qartod_time_flag:flag_values = "1, 2, 3, 4, 9" ;
		qartod_time_flag:ioos_category = "Other" ;
		qartod_time_flag:long_name = "" ;
		qartod_time_flag:standard_name = "" ;
	double semi_major_axis(obs) ;
		semi_major_axis:_FillValue = -9999.9 ;
		semi_major_axis:coordinates = "time z lon lat" ;
		semi_major_axis:long_name = "Error semi-major axis" ;
		semi_major_axis:units = "m" ;
		semi_major_axis:comment = "If the estimated position error is best expressed as an ellipse, this field gives the length in meters of the semi-major elliptical axis (one half of the major axis)." ;
		semi_major_axis:instrument = "instrument_location" ;
		semi_major_axis:platform = "platform" ;
	double semi_minor_axis(obs) ;
		semi_minor_axis:_FillValue = -9999.9 ;
		semi_minor_axis:coordinates = "time z lon lat" ;
		semi_minor_axis:long_name = "Error semi-minor axis" ;
		semi_minor_axis:units = "m" ;
		semi_minor_axis:comment = "If the estimated position error is best expressed as an ellipse, this field gives the length in meters of the semi-minor elliptical axis (one half of the minor axis)." ;
		semi_minor_axis:instrument = "instrument_location" ;
		semi_minor_axis:platform = "platform" ;
	double time(obs) ;
		time:_FillValue = -9999.9 ;
		time:units = "seconds since 1990-01-01 00:00:00Z" ;
		time:standard_name = "time" ;
		time:axis = "T" ;
		time:_CoordinateAxisType = "Time" ;
		time:calendar = "standard" ;
		time:ioos_category = "Time" ;
		time:long_name = "Time" ;
		time:actual_min = "2019-11-29T15:05:02Z" ;
		time:actual_max = "2020-04-27T08:29:22Z" ;
	int z(obs) ;
		z:_FillValue = -9999 ;
		z:axis = "Z" ;
		z:long_name = "depth" ;
		z:positive = "down" ;
		z:standard_name = "depth" ;
		z:units = "m" ;
		z:actual_min = 0. ;
		z:actual_max = 0. ;
		z:instrument = "instrument_location" ;
		z:platform = "platform" ;

// global attributes:
		:date_created = "2020-04-27T16:04:41Z" ;
		:featureType = "trajectory" ;
		:cdm_data_type = "Trajectory" ;
		:geospatial_bounds_vertical_crs = "EPSG:4326" ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_vertical_positive = "down" ;
		:naming_authority = "gov.noaa.ioos.atn" ;
		:publisher_email = "atndata@ioos.us" ;
		:publisher_name = "IOOS ATN" ;
		:publisher_url = "https://atn.ioos.us" ;
		:source = "Service Argos" ;
		:standard_name_vocabulary = "CF-v58" ;
		:geospatial_bbox = "POLYGON ((250.83 50.6209, 250.83 66.83069999999999, 159.0115000000001 66.83069999999999, 159.0115000000001 50.6209, 250.83 50.6209))" ;
		:geospatial_bounds = "POLYGON ((159.0115000000001 50.6209, 209.0858 59.7264, 250.83 66.83069999999999, 208.0173 58.7985, 160.9647 50.8049, 159.0115000000001 50.6209))" ;
		:geospatial_bounds_crs = "EPSG:4326" ;
		:geospatial_vertical_units = "m" ;
		:time_coverage_start = "2019-11-29T15:05:02Z" ;
		:time_coverage_end = "2020-04-27T08:29:22Z" ;
		:time_coverage_duration = "P149DT17H24M20S" ;
		:time_coverage_resolution = "P0DT0H42M21S" ;
		:date_issued = "2020-04-27T16:04:41Z" ;
		:date_modified = "2020-04-27T16:04:41Z" ;
		:argos_program_number = "11691" ;
		:creator_email = "michael.rehberg@alaska.gov" ;
		:first_uplink_date = "1575510820" ;
		:id = "5deb0b1d6321be14905284b8" ;
		:last_uplink_date = "1587997825" ;
		:ptt = "180473" ;
		:last_location_lat = "59.1356" ;
		:last_location_lon = "-151.4463" ;
		:last_location_date = "1587997825" ;
		:Conventions = "CF-1.6, ACDD-1.3" ;
		:acknowledgement = "NOAA IOOS, Axiom Data Science, Navy ONR,N OAA NMFS, Wildlife Computers, Argos" ;
		:creator_name = "Michael Rehberg" ;
		:creator_url = "https://www.adfg.alaska.gov/index.cfm?adfg=marinemammalprogram.stellerprogram" ;
		:infoUrl = "https://dev.axiomdatascience.com/?portal_id=99#search?type_group=all&query=habitat%20use%20of%20adult%20female%20steller&page=1" ;
		:institution = "Alaska Department of Fish and Game" ;
		:keywords = "atn,ioos,trajectory, steller sea lion" ;
		:license = "This animal telemery deployment data from Argos program 11691 and ptt 180473 is made available under the Open Database License: http://opendatacommons.org/licenses/odbl/1.0/. Any rights in individual contents of the database are licensed under the Database Contents License: http://opendatacommons.org/licenses/dbcl/1.0/" ;
		:metadata_link = "https://www.somelinkwhenwehaveacollectionpageat.NCEI.gov" ;
		:processing_level = "ATN DAC level 1 data prodcut [data levels yet to be explicitly documented[" ;
		:project = "Habitat Use of Adult Female Steller Sea Lions in the Endangered Western Distinct Population Segment, 2019-2020" ;
		:geospatial_lat_min = "50.6209" ;
		:geospatial_lat_max = "66.8307" ;
		:geospatial_lon_min = "-154.258" ;
		:geospatial_lon_max = "160.9647" ;
		:geospatial_vertical_min = "0.0" ;
		:geospatial_vertical_max = "0.0" ;
		:creator_country = "USA" ;
		:creator_institution = "Alaska Department of Fish and Game" ;
		:creator_sector = "gov_state" ;
		:date_metadata_modified = "2020-12-02T01:01:41Z" ;
		:instrument = "satellite telemetry tag" ;
		:platform = "animal" ;
		:platform_id = "5deb0b1d6321be14905284b8" ;
		:platform_name = "5deb0b1d6321be14905284b8" ;
		:platform_vocabulary = "https://mmisw.org/ont/ioos/platform" ;
		:program = "IOOS Animal Telemetry Network" ;
		:publisher_country = "USA" ;
		:publisher_institution = "US ATN DAC" ;
		:publisher_type = "institution" ;
		:vendor = "Wildlife Computers" ;
		:vendor_id = "5deb0b1d6321be14905284b8" ;
		:wmo_platform_code = "99nnnnn" ;
		:comment = "Flat Island, Alaska. Adult female with nursing pup (young-of-year). Brand X429. Mass not measured. \"SPLASH 10\" GPS location- and behavior-recording instrument glued to fur on top of the head." ;
		:sea_name = "North Pacific Ocean, Sea Okhotsk, and Bering Sea" ;
		:summary = "Wildlife Computers Splash 10 tag deployed on a Steller sea lion [Eumetopias jubatus] by Michael Rehberg in North Pacific Ocean, Sea Okhotsk, and Bering Sea from 2019-11-29 to 2020-04-27. PTT tag number 180473." ;
		:title = "Steller sea lion (Eumetopias jubatus) tag deployment from 2019-11-29 to 2020-04-27 in the North Pacific Ocean, Sea Okhotsk, and Bering Sea, ptt 180473" ;
		:history = "Mon Feb  8 14:31:10 2021: ncatted -a platform_groups,global,d,, Downloads/NCEI_test.2.nc Downloads/NCEI_test.3.nc\nMon Feb  8 14:28:47 2021: ncatted -a platform_category,global,d,, Downloads/NCEI_test.nc Downloads/NCEI_test.2.nc\nMon Feb  8 14:06:17 2021: ncks -x -v instrument,trajectory,deploy_id,type,comment,qartod_rollup_flag Downloads/atn_deployment_01.5.nc Downloads/atn_deployment_NCEI_test.nc\nnarrative description of ATN DAC processes for creating this file and sending to NCEI" ;
		:NCO = "4.7.2" ;
}