netcdf ATN_Trajectory {
dimensions:
	obs = < dim1 > ; //..........................................................................Total number of observations
	strlen_taxon_name = < dim2 > ; //............................................................Length of the taxon name string (eg. 18 for "Eumetopias jubatus")
	strlen_taxon_lsid = < dim3 > ; //............................................................Length of the taxon lsid string (eg. 41 for "urn:lsid:marinespecies.org:taxname:254999")
variables:
	double time(obs) ;
		time:_FillValue = "" ;
		time:units = "" ;
		time:standard_name = "" ;
		time:axis = "" ;
		time:_CoordinateAxisType = "" ;
		time:calendar = "" ;
		time:ioos_category = "" ;
		time:long_name = "" ;
		time:actual_min = "" ;
		time:actual_max = "" ;
	int z(obs) ;
		zi:_FillValue = "" ;
		z:axis = "" ;
		z:long_name = "" ;
		z:positive = "" ;
		z:standard_name = "" ;
		z:units = "" ;
		z:actual_min = "" ;
		z:actual_max = "" ;
		z:instrument = "instrument_pressure" ;
		z:platform = "animal" ;
	double lat(obs) ;
		lat:_FillValue = "" ;
		lat:axis = "" ;
		lat:_CoordinateAxisType = "" ;
		lat:ioos_category = "" ;
		lat:long_name = "" ;
		lat:standard_name = "" ;
		lat:units = "" ;
		lat:valid_max = "" ;
		lat:valid_min = "" ;
		lat:actual_min = "" ;
		lat:actual_max = "" ;
		lat:instrument = "instrument_location" ;
		lat:platform = "animal" ;
	double lon(obs) ;
		lon:_FillValue = "" ;
		lon:axis = "" ;
		lon:_CoordinateAxisType = "" ;
		lon:ioos_category = "" ;
		lon:long_name = "" ;
		lon:standard_name = "" ;
		lon:units = "" ;
		lon:valid_max = "" ;
		lon:valid_min = "" ;
		lon:actual_min = "" ;
		lon:actual_max = "" ;
		lon:instrument = "instrument_location" ;
		lon:platform = "animal" ;
	string location_class(obs) ;
		location_class:coordinates = "" ;
		location_class:long_name = "" ;
		location_class:standard_name = "" ;
		location_class:ioos_category = "" ;
		location_class:comment = "" ;
		location_class:code_values = "" ;
		location_class:code_meanings = "" ;
		location_class:instrument = "instrument_location" ;
		location_class:platform = "animal" ;
	string instrument_tag ;
		instrument_tag:long_name = "" ;
		instrument_tag:comment = "" ;
		instrument_tag:manufacturer = "" ;
		instrument_tag:make_model = "" ;
		instrument_tag:calibration_date = "" ;
		instrument_tag:serial_number = "" ;
	string instrument_location ;
		instrument_location:long_name = "" ;
		instrument_location:location_type = "" ;
		instrument_location:comment = "" ;
		instrument_location:manufacturer = "" ;
		instrument_location:make_model = "" ;
		instrument_location:calibration_date = "" ;
		instrument_location:serial_number = "" ;
	string instrument_pressure ;
		instrument_pressure:long_name = "" ;
		instrument_pressure:comment = "" ;
		instrument_pressure:manufacturer = "" ;
		instrument_pressure:make_model = "" ;
		instrument_pressure:calibration_date = "" ;
		instrument_pressure:serial_number = "" ;
	string animal ; //.........................................................................Treated as a platform container variable
		animal:cf_role = "" ;
		animal:long_name = "" ;
		animal:platform_type = "" ;
		animal:platform_vocabulary = "" ;
		animal:valid_name = "" ;
		animal:AphiaID = "" ;
		animal:scientificname = "" ;
		animal:authority = "" ;
		animal:kingdom = "" ;
		animal:phylum = "" ;
		animal:class = "" ;
		animal:order = "" ;
		animal:family = "" ;
		animal:genus = "" ;
		animal:rank = "" ;
		animal:superdomain = "" ;
		animal:subphylum = "" ;
		animal:superclass = "" ;
		animal:subclass = "" ;
		animal:suborder = "" ;
		animal:infraorder = "" ;
		animal:species = "" ;
		animal:taxonRankID = "" ;
	string taxon_name(strlen_taxon_name) ;  //.................................................Eg. "Eumetopias jubatus"
	    	taxon_name:standard_name = "biological_taxon_name" ;
	    	taxon_name:long_name = "" ; //.....................................................most precise taxonomic classification
	string taxon_lsid(strlen_taxon_lsid) ;  //.................................................Eg. "urn:lsid:marinespecies.org:taxname:254999"
	    	taxon_lsid:standard_name = "biological_taxon_id" ;
	    	taxon_lsid:long_name = "Taxon identifier" ;
	    	taxon_lsid:source = "" ; //........................................................source of the lsid (eg. WoRMS, ITIS)
	double ellipse_orientation(obs) ;
		ellipse_orientation:_FillValue = "" ;
		ellipse_orientation:coordinates = "" ;
		ellipse_orientation:long_name = "" ;
		ellipse_orientation:units = "" ;
		ellipse_orientation:comment = "" ;
		ellipse_orientation:instrument = "" ;
		ellipse_orientation:platform = "animal" ;
	double error_radius(obs) ;
		error_radius:_FillValue = "" ;
		error_radius:coordinates = "" ;
		error_radius:long_name = "" ;
		error_radius:units = "" ;
		error_radius:comment = "" ;
		error_radius:instrument = "" ;
		error_radius:platform = "animal" ;
	double semi_major_axis(obs) ;
		semi_major_axis:_FillValue = "" ;
		semi_major_axis:coordinates = "" ;
		semi_major_axis:long_name = "" ;
		semi_major_axis:units = "" ;
		semi_major_axis:comment = "" ;
		semi_major_axis:instrument = "instrument_location" ;
		semi_major_axis:platform = "animal" ;
	double semi_minor_axis(obs) ;
		semi_minor_axis:_FillValue = "" ;
		semi_minor_axis:coordinates = "" ;
		semi_minor_axis:long_name = "" ;
		semi_minor_axis:units = "" ;
		semi_minor_axis:comment = "" ;
		semi_minor_axis:instrument = "instrument_location" ;
		semi_minor_axis:platform = "animal" ;
	double offset(obs) ;
		offset:_FillValue = "" ;
		offset:coordinates = "" ;
		offset:long_name = "" ;
		offset:units = "" ;
		offset:comment = "" ;
	double offset_orientation(obs) ;
		offset_orientation:_FillValue = "" ;
		offset_orientation:coordinates = "" ;
		offset_orientation:long_name = "" ;
		offset_orientation:units = "" ;
		offset_orientation:comment = "" ;
	int crs ;
		crs:epsg_code = "" ;
		crs:grid_mapping_name = "" ;
		crs:inverse_flattening = "" ;
		crs:ioos_category = "" ;
		crs:long_name = "" ;
		crs:semi_major_axis = "" ;
	string qartod_rollup_flag(obs) ;
		qartod_rollup_flag:_FillValue = "" ;
		qartod_rollup_flag:flag_meanings = "" ;
		qartod_rollup_flag:flag_values = "" ;
		qartod_rollup_flag:ioos_category = "" ;
		qartod_rollup_flag:long_name = "" ;
		qartod_rollup_flag:standard_name = "" ;
	string qartod_speed_flag(obs) ;
		qartod_speed_flag:_FillValue = "" ;
		qartod_speed_flag:flag_meanings = "" ;
		qartod_speed_flag:flag_values = "" ;
		qartod_speed_flag:ioos_category = "" ;
		qartod_speed_flag:long_name = "" ;
		qartod_speed_flag:standard_name = "" ;
	string qartod_location_flag(obs) ;
		qartod_location_flag:_FillValue = "" ;
		qartod_location_flag:flag_meanings = "" ;
		qartod_location_flag:flag_values = "" ;
		qartod_location_flag:ioos_category = "" ;
		qartod_location_flag:long_name = "" ;
		qartod_location_flag:standard_name = "" ;
	string qartod_time_flag(obs) ;
		qartod_time_flag:_FillValue = "" ;
		qartod_time_flag:flag_meanings = "" ;
		qartod_time_flag:flag_values = "" ;
		qartod_time_flag:ioos_category = "" ;
		qartod_time_flag:long_name = "" ;
		qartod_time_flag:standard_name = "" ;

// global attributes:
		:argos_program_number = "" ;
		:acknowledgement = "" ;
		:cdm_data_type = "" ;
		:comment = "" ;
		:common_name = "" ;
		:Conventions = "" ;
		:creator_country = "" ;
		:creator_email = "" ;
		:creator_institution = "" ;
		:creator_name = "" ;
		:creator_sector = "" ;
		:creator_url = "" ;
		:date_created = "" ;
		:date_issued = "" ;
		:date_modified = "" ;
		:date_metadata_modified = "" ;
		:featureType = "" ;
		:first_uplink_date = "" ;
		:geospatial_bbox = "" ;
		:geospatial_bounds_vertical_crs = "" ;
		:geospatial_lat_units = "" ;
		:geospatial_lon_units = "" ;
		:geospatial_vertical_positive = "" ;
		:geospatial_bounds = "" ;
		:geospatial_bounds_crs = "" ;
		:geospatial_vertical_units = "" ;
		:geospatial_lat_min = "" ;
		:geospatial_lat_max = "" ;
		:geospatial_lon_min = "" ;
		:geospatial_lon_max = "" ;
		:geospatial_vertical_min = "" ;
		:geospatial_vertical_max = "" ;
		:history = "" ;
		:id = "" ;
		:infoUrl = "" ;
		:institution = "" ;
		:instrument = "" ;
		:keywords = "" ;
		:keywords_vocabulary = "" ;
		:naming_authority = "" ;
		:publisher_email = "" ;
		:publisher_name = "" ;
		:publisher_url = "" ;
		:source = "" ;
		:standard_name_vocabulary = "" ;
		:time_coverage_start = "" ;
		:time_coverage_end = "" ;
		:time_coverage_duration = "" ;
		:time_coverage_resolution = "" ;
		:last_uplink_date = "" ;
		:last_location_lat = "" ;
		:last_location_lon = "" ;
		:last_location_date = "" ;
		:license = "" ;
		:metadata_link = "" ;
		:NCO = "" ;
		:processing_level = "" ;
		:project = "" ;
		:platform = "animal" ;
		:platform_id = "" ;
		:platform_name = "" ;
		:platform_vocabulary = "" ;
		:program = "" ;
		:ptt = "" ;
		:publisher_country = "" ;
		:publisher_institution = "" ;
		:publisher_type = "" ;
		:sea_name = "" ;
		:summary = "" ;
		:title = "" ;
		:vendor = "" ;
		:vendor_id = "" ;
		:wmo_platform_code = "" ;
		
}
