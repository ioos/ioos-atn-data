netcdf atn_trajectory_template {
dimensions:
	time = 1 ; //..........................................................................Total number of observations
	strlen_taxon_name = 1 ; //............................................................Length of the taxon name string (eg. 18 for "Eumetopias jubatus")
	strlen_taxon_lsid = 1 ; //............................................................Length of the taxon lsid string (eg. 41 for "urn:lsid:marinespecies.org:taxname:254999")
variables:
	string trajectory ;
		trajectory:cf_role = "trajectory_id" ;
		trajectory:long_name = "trajectory identifier" ;
	double time(time) ;
		time:_FillValue = -9999.9 ;
		time:units = "seconds since 1990-01-01 00:00:00Z" ;
		time:standard_name = "time" ;
		time:axis = "T" ;
		time:_CoordinateAxisType = "Time" ;
		time:calendar = "" ;
		time:long_name = "Time" ;
		time:actual_min = "" ;
		time:actual_max = "" ;
		time:ancillary_variables = "qartod_time_flag qartod_rollup_flag" ;
	int z(time) ;
		z:_FillValue = -9999 ;
		z:axis = "Z" ;
		z:long_name = "depth" ;
		z:positive = "down" ;
		z:standard_name = "depth" ;
		z:units = "m" ;
		z:actual_min = "" ;
		z:actual_max = "" ;
		z:instrument = "instrument_pressure" ;
		z:platform = "animal" ;
	double lat(time) ;
		lat:_FillValue = -9999 ;
		lat:axis = "Y" ;
		lat:_CoordinateAxisType = "Lat" ;
		lat:long_name = "Profile location latitude" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:valid_max = 90. ;
		lat:valid_min = -90. ;
		lat:actual_min = "" ;
		lat:actual_max = "" ;
		lat:instrument = "instrument_location" ;
		lat:platform = "animal" ;
		lat:ancillary_variables = "qartod_location_flag qartod_rollup_flag" ;
	double lon(time) ;
		lon:_FillValue = -9999 ;
		lon:axis = "X" ;
		lon:_CoordinateAxisType = "Lon" ;
		lon:long_name = "Profile location longitude" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:valid_max = 180. ;
		lon:valid_min = -180. ;
		lon:actual_min = "" ;
		lon:actual_max = "" ;
		lon:instrument = "instrument_location" ;
		lon:platform = "animal" ;
		lon:ancillary_variables = "qartod_location_flag qartod_rollup_flag" ;
	string location_class(time) ;
		location_class:coordinates = "time z lon lat" ;
		location_class:long_name = "Location Quality Code" ;
		location_class:standard_name = "status_flag" ;
		location_class:comment = "Quality codes from the ARGOS satellite (in meters): G,3,2,1,0,A,B,Z. See http://www.argos-system.org/manual/3-location/34_location_classes.htm" ;
		location_class:code_values = "G,3,2,1,0,A,B,Z" ;
		location_class:code_meanings = "estimated error less than 100m and 1+ messages received per satellite pass,estimated error less than 250m and 4+ messages received per satellite pass,estimated error between 250m and 500m and 4+ messages per satellite pass,estimated error between 500m and 1500m and 4+ messages per satellite pass,estimated error greater than 1500m and 4+ messages received per satellite pass,no least squares estimated error or unbounded kalman filter estimated error and 3 messages received per satellite pass,no least squares estimated error or unbounded kalman filter estimated error and 1 or 2 messages received per satellite pass,invalid location (available for Service Plus or Auxilliary Location Processing)" ;
		location_class:instrument = "instrument_location" ;
		location_class:platform = "animal" ;
		location_class:ancillary_variables = "qartod_location_flag qartod_rollup_flag" ;
	double ellipse_orientation(time) ;
		ellipse_orientation:_FillValue = -9999.9 ;
		ellipse_orientation:coordinates = "time z lon lat" ;
		ellipse_orientation:long_name = "Ellipse orientation" ;
		ellipse_orientation:units = "degrees" ;
		ellipse_orientation:comment = "The angle in degrees of the ellipse from true north, proceeding clockwise (0 to 360). A blank field represents 0 degrees." ;
		ellipse_orientation:instrument = "instrument_location" ;
		ellipse_orientation:platform = "animal" ;
	double error_radius(time) ;
		error_radius:_FillValue = -9999.9 ;
		error_radius:coordinates = "time z lon lat" ;
		error_radius:long_name = "Error radius" ;
		error_radius:units = "m" ;
		error_radius:comment = "If the position is best represented as a circle, this field gives the radius of that circle in meters." ;
		error_radius:instrument = "instrument_location" ;
		error_radius:platform = "animal" ;
	double semi_major_axis(time) ;
		semi_major_axis:_FillValue = -9999.9 ;
		semi_major_axis:coordinates = "time z lon lat" ;
		semi_major_axis:long_name = "Error semi-major axis" ;
		semi_major_axis:units = "m" ;
		semi_major_axis:comment = "If the estimated position error is best expressed as an ellipse, this field gives the length in meters of the semi-major elliptical axis (one half of the major axis)." ;
		semi_major_axis:instrument = "instrument_location" ;
		semi_major_axis:platform = "animal" ;
	double semi_minor_axis(time) ;
		semi_minor_axis:_FillValue = -9999.9 ;
		semi_minor_axis:coordinates = "time z lon lat" ;
		semi_minor_axis:long_name = "Error semi-minor axis" ;
		semi_minor_axis:units = "m" ;
		semi_minor_axis:comment = "If the estimated position error is best expressed as an ellipse, this field gives the length in meters of the semi-minor elliptical axis (one half of the minor axis)." ;
		semi_minor_axis:instrument = "instrument_location" ;
		semi_minor_axis:platform = "animal" ;
	double offset(time) ;
		offset:_FillValue = -9999.9 ;
		offset:coordinates = "time z lon lat" ;
		offset:long_name = "Offset" ;
		offset:units = "m" ;
		offset:comment = "This field is non-zero if the circle or ellipse are not centered on the (Latitude, Longitude) values on this row. \"Offset\" gives the distance in meters from (Latitude, Longitude) to the center of the ellipse." ;
		offset:instrument = "instrument_location" ;
		offset:platform = "platform" ;
	double offset_orientation(time) ;
		offset_orientation:_FillValue = -9999.9 ;
		offset_orientation:coordinates = "time z lon lat" ;
		offset_orientation:long_name = "Offset orientation" ;
		offset_orientation:units = "degrees" ;
		offset_orientation:comment = "If the \"Offset\" field is non-zero, this field is the angle in degrees from (Latitude, Longitude) to the center of the ellipse. Zero degrees is true north; a blank field represents 0 degrees." ;
		offset_orientation:instrument = "instrument_location" ;
		offset_orientation:platform = "platform" ;
	int64 qartod_rollup_flag(time) ;
		qartod_rollup_flag:_FillValue = "" ;
		qartod_rollup_flag:flag_meanings = "PASS NOT_EVALUATED SUSPECT FAIL MISSING" ;
		qartod_rollup_flag:flag_values = "1, 2, 3, 4, 9" ;
		qartod_rollup_flag:long_name = "" ;
		qartod_rollup_flag:standard_name = "aggregate_quality_flag" ;
		qartod_rollup_flag:references = "" ;
	int64 qartod_speed_flag(time) ;
		qartod_speed_flag:_FillValue = "" ;
		qartod_speed_flag:flag_meanings = "PASS NOT_EVALUATED SUSPECT FAIL MISSING" ;
		qartod_speed_flag:flag_values = "1, 2, 3, 4, 9" ;
		qartod_speed_flag:long_name = "" ;
		qartod_speed_flag:standard_name = "gross_range_test_quality_flag" ;
		qartod_speed_flag:references = "" ;
	int64 qartod_location_flag(time) ;
		qartod_location_flag:_FillValue = "" ;
		qartod_location_flag:flag_meanings = "PASS NOT_EVALUATED SUSPECT FAIL MISSING" ;
		qartod_location_flag:flag_values = "1, 2, 3, 4, 9" ;
		qartod_location_flag:long_name = "" ;
		qartod_location_flag:standard_name = "location_test_quality_flag" ;
		qartod_location_flag:references = "" ;
	int64 qartod_time_flag(time) ;
		qartod_time_flag:_FillValue = "" ;
		qartod_time_flag:flag_meanings = "PASS NOT_EVALUATED SUSPECT FAIL MISSING" ;
		qartod_time_flag:flag_values = "1, 2, 3, 4, 9" ;
		qartod_time_flag:long_name = "" ;
		qartod_time_flag:standard_name = "gross_range_test_quality_flag" ;
		qartod_time_flag:references = "" ;
	string taxon_name(strlen_taxon_name) ;  //.................................................Eg. "Eumetopias jubatus"
	    taxon_name:standard_name = "biological_taxon_name" ;
	    taxon_name:long_name = "" ; //.....................................................most precise taxonomic classification
	string taxon_lsid(strlen_taxon_lsid) ;  //.................................................Eg. "urn:lsid:marinespecies.org:taxname:254999"
	    taxon_lsid:standard_name = "biological_taxon_lsid" ;//.............................CF table 76/77 incorrectly lists this as biological_taxon_identifier
	    taxon_lsid:long_name = "Taxon identifier" ;
	    taxon_lsid:source = "" ; //........................................................source of the lsid (eg. WoRMS, ITIS)
	string instrument_tag ;
		instrument_tag:long_name = "" ;
		instrument_tag:comment = "" ;
		instrument_tag:manufacturer = "" ;
		instrument_tag:make_model = "" ;
		instrument_tag:calibration_date = "" ;
		instrument_tag:serial_number = "" ;
	string instrument_location ;
		instrument_location:long_name = "" ;
		instrument_location:location_type = "" ;
		instrument_location:comment = "" ;
		instrument_location:manufacturer = "" ;
		instrument_location:make_model = "" ;
		instrument_location:calibration_date = "" ;
		instrument_location:serial_number = "" ;
	string instrument_pressure ;
		instrument_pressure:long_name = "" ;
		instrument_pressure:comment = "" ;
		instrument_pressure:manufacturer = "" ;
		instrument_pressure:make_model = "" ;
		instrument_pressure:calibration_date = "" ;
		instrument_pressure:serial_number = "" ;
	string animal ; //.........................................................................Treated as a platform container variable
		animal:long_name = "" ;
		animal:valid_name = "" ;
		animal:AphiaID = "" ;
		animal:scientificname = "" ;
		animal:authority = "" ;
		animal:kingdom = "" ;
		animal:phylum = "" ;
		animal:class = "" ;
		animal:order = "" ;
		animal:family = "" ;
		animal:genus = "" ;
		animal:rank = "" ;
		animal:superdomain = "" ;
		animal:subphylum = "" ;
		animal:superclass = "" ;
		animal:subclass = "" ;
		animal:suborder = "" ;
		animal:infraorder = "" ;
		animal:species = "" ;
		animal:taxonRankID = "" ;
	int crs ;
		crs:epsg_code = "EPSG:4326" ;
		crs:grid_mapping_name = "latitude_longitude" ;
		crs:inverse_flattening = 298.257223563 ;
		crs:ioos_category = "Other" ;
		crs:long_name = "http://www.opengis.net/def/crs/EPSG/0/4326" ;
		crs:semi_major_axis = 6378137. ;

// global attributes:
		:argos_program_number = "" ;
		:acknowledgement = "" ;
		:cdm_data_type = "Trajectory" ;
		:comment = "" ;
		:common_name = "" ;
		:Conventions = "CF-1.6, ACDD-1.3, IOOS-1.2" ;
		:creator_country = "" ;
		:creator_email = "" ;
		:creator_institution = "" ;
		:creator_name = "" ;
		:creator_sector = "" ;
		:creator_url = "" ;
		:date_created = "" ;
		:date_issued = "" ;
		:date_modified = "" ;
		:date_metadata_modified = "" ;
		:featureType = "trajectory" ;
		:first_uplink_date = "" ;
		:geospatial_bbox = "" ;
		:geospatial_bounds_vertical_crs = "" ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_vertical_positive = "down" ;
		:geospatial_bounds = "" ;
		:geospatial_bounds_crs = "" ;
		:geospatial_vertical_units = "m" ;
		:geospatial_lat_min = "" ;
		:geospatial_lat_max = "" ;
		:geospatial_lon_min = "" ;
		:geospatial_lon_max = "" ;
		:geospatial_vertical_min = "" ;
		:geospatial_vertical_max = "" ;
		:history = "" ;
		:id = "" ;
		:infoUrl = "" ;
		:institution = "" ;
		:instrument = "" ;
		:keywords = "EARTH SCIENCE > BIOLOGICAL CLASSIFICATION > ANIMALS/INVERTEBRATES" ;
		:keywords_vocabulary = "GCMD Earth Science Keywords. Version 10.0" ;
		:naming_authority = "" ;
		:ncei_template_version = "NCEI_NetCDF_Trajectory_Template_v2.0" ;
		:publisher_email = "" ;
		:publisher_name = "" ;
		:publisher_url = "" ;
		:source = "" ;
		:standard_name_vocabulary = "CF Standard Name Table v77" ;
		:time_coverage_start = "" ;
		:time_coverage_end = "" ;
		:time_coverage_duration = "" ;
		:time_coverage_resolution = "" ;
		:last_uplink_date = "" ;
		:last_location_lat = "" ;
		:last_location_lon = "" ;
		:last_location_date = "" ;
		:license = "" ;
		:metadata_link = "" ;
		:NCO = "" ;
		:processing_level = "" ;
		:project = "" ;
		:platform = "animal" ;
		:platform_id = "" ;
		:platform_name = "" ;
		:platform_vocabulary = "" ;
		:program = "" ;
		:ptt = "" ;
		:publisher_country = "" ;
		:publisher_institution = "" ;
		:publisher_type = "" ;
		:sea_name = "" ;
		:summary = "This is a template file for the IOOS Animal Telemetry Network (ATN) trajectory observations." ;
		:title = "Animal Telemetry Network trajectory netCDF file template" ;
		:vendor = "" ;
		:vendor_id = "" ;
		:wmo_platform_code = "" ;
		
}
